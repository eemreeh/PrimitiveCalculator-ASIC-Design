* NGSPICE file created from PrimitiveCalculator.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtn_1 abstract view
.subckt sky130_fd_sc_hd__dlxtn_1 D GATE_N VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtn_2 abstract view
.subckt sky130_fd_sc_hd__dlxtn_2 D GATE_N VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtp_1 abstract view
.subckt sky130_fd_sc_hd__dlxtp_1 D GATE VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

.subckt PrimitiveCalculator VGND VPWR clk led_flag restart rotary_a rotary_b rst select
+ seven_segment_digit seven_segment_out[0] seven_segment_out[1] seven_segment_out[2]
+ seven_segment_out[3] seven_segment_out[4] seven_segment_out[5] seven_segment_out[6]
XFILLER_36_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1270_ _1270_/A _1270_/B VGND VGND VPWR VPWR _1271_/B sky130_fd_sc_hd__and2_1
XFILLER_51_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0985_ _0985_/A _0985_/B VGND VGND VPWR VPWR _1028_/A sky130_fd_sc_hd__nor2_1
X_1606_ _1603_/A _1588_/X _1605_/Y _1599_/X VGND VGND VPWR VPWR _1768_/D sky130_fd_sc_hd__o211a_1
X_1399_ _1399_/A _1399_/B VGND VGND VPWR VPWR _1400_/B sky130_fd_sc_hd__nor2_1
X_1468_ _1516_/A _1523_/A _1538_/B VGND VGND VPWR VPWR _1468_/X sky130_fd_sc_hd__a21o_1
X_1537_ _1537_/A VGND VGND VPWR VPWR _1820_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_63_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1253_ _1821_/Q _1282_/B _1253_/C VGND VGND VPWR VPWR _1253_/X sky130_fd_sc_hd__and3_1
X_1322_ _1426_/C _1323_/B _1446_/B VGND VGND VPWR VPWR _1322_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_64_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1184_ _1202_/A _1184_/B _1195_/A VGND VGND VPWR VPWR _1184_/X sky130_fd_sc_hd__and3b_1
XFILLER_17_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0968_ _0968_/A _0968_/B _0968_/C _0968_/D VGND VGND VPWR VPWR _1004_/A sky130_fd_sc_hd__or4_1
XFILLER_32_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0899_ _1830_/Q _1831_/Q VGND VGND VPWR VPWR _0921_/B sky130_fd_sc_hd__nor2_1
XFILLER_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1305_ _1821_/Q _1282_/B _1348_/D _1388_/B VGND VGND VPWR VPWR _1305_/X sky130_fd_sc_hd__a22o_1
XFILLER_37_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1236_ _1246_/B _1263_/B VGND VGND VPWR VPWR _1238_/A sky130_fd_sc_hd__nor2_1
X_1098_ _1142_/A _1142_/B _1098_/C _1098_/D VGND VGND VPWR VPWR _1100_/A sky130_fd_sc_hd__or4_1
X_1167_ input4/X VGND VGND VPWR VPWR _1727_/B sky130_fd_sc_hd__inv_2
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1021_ _1057_/A _1057_/B _1392_/B VGND VGND VPWR VPWR _1059_/B sky130_fd_sc_hd__a21o_1
XFILLER_34_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1785_ _1839_/CLK _1785_/D VGND VGND VPWR VPWR _1785_/Q sky130_fd_sc_hd__dfxtp_1
X_1854_ _1816_/Q _1854_/D VGND VGND VPWR VPWR _1854_/Q sky130_fd_sc_hd__dfxtp_1
X_1219_ _1388_/B VGND VGND VPWR VPWR _1426_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_44_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1570_ _1570_/A VGND VGND VPWR VPWR _1760_/D sky130_fd_sc_hd__clkbuf_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1004_ _1004_/A _1004_/B VGND VGND VPWR VPWR _1006_/B sky130_fd_sc_hd__and2_1
X_1837_ _1837_/CLK _1837_/D VGND VGND VPWR VPWR _1837_/Q sky130_fd_sc_hd__dfxtp_1
X_1768_ _1816_/Q _1768_/D VGND VGND VPWR VPWR _1768_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1699_ _1697_/X _1698_/X _1803_/Q _1456_/A VGND VGND VPWR VPWR _1699_/X sky130_fd_sc_hd__o211a_1
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput7 _1835_/Q VGND VGND VPWR VPWR seven_segment_digit sky130_fd_sc_hd__buf_2
XFILLER_63_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1622_ _1619_/X _1620_/X _1621_/Y VGND VGND VPWR VPWR _1622_/X sky130_fd_sc_hd__a21o_1
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1553_ _1553_/A VGND VGND VPWR VPWR _1804_/D sky130_fd_sc_hd__clkbuf_1
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1484_ _1512_/B VGND VGND VPWR VPWR _1505_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_54_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0984_ _1244_/A _0983_/X _0947_/Y VGND VGND VPWR VPWR _0985_/B sky130_fd_sc_hd__a21o_1
X_1605_ _1628_/A _1605_/B VGND VGND VPWR VPWR _1605_/Y sky130_fd_sc_hd__nand2_1
X_1536_ _1536_/A _1538_/B VGND VGND VPWR VPWR _1537_/A sky130_fd_sc_hd__and2_1
X_1398_ _1398_/A _1398_/B _1398_/C VGND VGND VPWR VPWR _1399_/B sky130_fd_sc_hd__nor3_1
X_1467_ _1540_/A VGND VGND VPWR VPWR _1538_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1252_ _1388_/B _1304_/B VGND VGND VPWR VPWR _1255_/A sky130_fd_sc_hd__nand2_1
X_1321_ _1210_/X _1293_/Y _1294_/X _1320_/X _1195_/X VGND VGND VPWR VPWR _1321_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1183_ _1183_/A _1806_/Q VGND VGND VPWR VPWR _1195_/A sky130_fd_sc_hd__nor2_1
X_0967_ _1162_/A _1823_/Q VGND VGND VPWR VPWR _0968_/D sky130_fd_sc_hd__and2_1
XFILLER_32_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0898_ _1833_/Q _1832_/Q _1834_/Q VGND VGND VPWR VPWR _0921_/A sky130_fd_sc_hd__nor3_2
X_1519_ _1536_/A _1532_/B _1523_/A VGND VGND VPWR VPWR _1520_/A sky130_fd_sc_hd__and3_1
XFILLER_55_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1304_ _1347_/A _1304_/B VGND VGND VPWR VPWR _1346_/A sky130_fd_sc_hd__nand2_1
XFILLER_37_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1235_ _1235_/A _1235_/B VGND VGND VPWR VPWR _1263_/B sky130_fd_sc_hd__nor2_1
X_1166_ _1161_/X _1163_/Y _1708_/A VGND VGND VPWR VPWR _1786_/D sky130_fd_sc_hd__a21oi_1
X_1097_ _1146_/A _1146_/B _1411_/B VGND VGND VPWR VPWR _1098_/D sky130_fd_sc_hd__a21oi_1
XFILLER_52_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1020_ _1020_/A VGND VGND VPWR VPWR _1392_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_42_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1784_ _1837_/CLK _1784_/D VGND VGND VPWR VPWR _1784_/Q sky130_fd_sc_hd__dfxtp_1
X_1853_ _1816_/Q _1853_/D VGND VGND VPWR VPWR _1853_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1149_ _1146_/Y _1148_/Y _1149_/S VGND VGND VPWR VPWR _1149_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1218_ _1193_/X _1194_/X _1211_/X _1214_/Y _1217_/X VGND VGND VPWR VPWR _1788_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1003_ _1348_/D VGND VGND VPWR VPWR _1221_/B sky130_fd_sc_hd__buf_2
X_1767_ _1816_/Q _1767_/D VGND VGND VPWR VPWR _1807_/D sky130_fd_sc_hd__dfxtp_2
X_1836_ _1837_/CLK _1836_/D VGND VGND VPWR VPWR _1836_/Q sky130_fd_sc_hd__dfxtp_1
X_1698_ _1854_/Q _1855_/Q _1856_/Q _1857_/Q VGND VGND VPWR VPWR _1698_/X sky130_fd_sc_hd__or4_1
XFILLER_57_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput10 _1506_/X VGND VGND VPWR VPWR seven_segment_out[2] sky130_fd_sc_hd__buf_2
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput8 _1497_/X VGND VGND VPWR VPWR seven_segment_out[0] sky130_fd_sc_hd__buf_2
XFILLER_63_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1552_ _1554_/A _1794_/Q _1556_/A VGND VGND VPWR VPWR _1553_/A sky130_fd_sc_hd__and3_1
X_1621_ _1619_/X _1620_/X _1596_/A VGND VGND VPWR VPWR _1621_/Y sky130_fd_sc_hd__o21ai_1
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1483_ _1777_/Q _1708_/B _1482_/X VGND VGND VPWR VPWR _1512_/B sky130_fd_sc_hd__o21a_1
X_1819_ _1819_/D _0880_/X VGND VGND VPWR VPWR _1819_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_45_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0983_ _1348_/C _0983_/B _0983_/C VGND VGND VPWR VPWR _0983_/X sky130_fd_sc_hd__or3_1
X_1604_ _1604_/A _1604_/B VGND VGND VPWR VPWR _1605_/B sky130_fd_sc_hd__xnor2_1
X_1535_ _1535_/A VGND VGND VPWR VPWR _1819_/D sky130_fd_sc_hd__clkbuf_1
X_1397_ _1398_/A _1398_/B _1398_/C VGND VGND VPWR VPWR _1399_/A sky130_fd_sc_hd__o21a_1
X_1466_ _1668_/B _1516_/A _1665_/A VGND VGND VPWR VPWR _1540_/A sky130_fd_sc_hd__nor3b_1
XFILLER_50_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1320_ _1320_/A _1320_/B VGND VGND VPWR VPWR _1320_/X sky130_fd_sc_hd__xor2_1
XFILLER_49_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1182_ _1158_/A _1421_/A _1137_/A _1382_/A VGND VGND VPWR VPWR _1184_/B sky130_fd_sc_hd__a22o_1
X_1251_ _1181_/A _1295_/A _1250_/X VGND VGND VPWR VPWR _1260_/A sky130_fd_sc_hd__o21ai_1
X_0966_ _0966_/A VGND VGND VPWR VPWR _1162_/A sky130_fd_sc_hd__buf_2
X_0897_ _1825_/Q VGND VGND VPWR VPWR _1327_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_59_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1449_ _1270_/A _1270_/B _1291_/B _1329_/A _1289_/A VGND VGND VPWR VPWR _1449_/X
+ sky130_fd_sc_hd__o311a_1
X_1518_ _1518_/A VGND VGND VPWR VPWR _1827_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1303_ _1426_/A _1198_/B _1255_/B _1253_/X VGND VGND VPWR VPWR _1338_/A sky130_fd_sc_hd__a31oi_2
X_1096_ _1411_/B _1146_/A _1146_/B VGND VGND VPWR VPWR _1098_/C sky130_fd_sc_hd__and3_1
XFILLER_37_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1234_ _1235_/A _1235_/B VGND VGND VPWR VPWR _1246_/B sky130_fd_sc_hd__and2_1
X_1165_ _1711_/S VGND VGND VPWR VPWR _1708_/A sky130_fd_sc_hd__clkbuf_2
X_0949_ _0962_/B _0949_/B VGND VGND VPWR VPWR _0953_/A sky130_fd_sc_hd__and2_1
XFILLER_43_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1852_ _1816_/Q _1852_/D VGND VGND VPWR VPWR _1852_/Q sky130_fd_sc_hd__dfxtp_1
X_1783_ _1837_/CLK _1783_/D VGND VGND VPWR VPWR _1783_/Q sky130_fd_sc_hd__dfxtp_1
X_1148_ _1098_/C _1098_/D _1147_/Y _1142_/A VGND VGND VPWR VPWR _1148_/Y sky130_fd_sc_hd__o22ai_1
X_1079_ _1205_/B _1114_/B _1122_/B _1133_/A _1078_/X VGND VGND VPWR VPWR _1082_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_52_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1217_ _1456_/A VGND VGND VPWR VPWR _1217_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_28_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1002_ _1112_/A _1024_/B VGND VGND VPWR VPWR _1039_/A sky130_fd_sc_hd__nand2_1
XFILLER_30_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1835_ _1816_/Q _1835_/D VGND VGND VPWR VPWR _1835_/Q sky130_fd_sc_hd__dfxtp_2
X_1766_ _1816_/Q _1766_/D VGND VGND VPWR VPWR _1806_/D sky130_fd_sc_hd__dfxtp_1
X_1697_ _1850_/Q _1851_/Q _1852_/Q _1853_/Q VGND VGND VPWR VPWR _1697_/X sky130_fd_sc_hd__or4_1
XFILLER_57_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput9 _1502_/Y VGND VGND VPWR VPWR seven_segment_out[1] sky130_fd_sc_hd__buf_2
Xoutput11 _1508_/Y VGND VGND VPWR VPWR seven_segment_out[3] sky130_fd_sc_hd__buf_2
XFILLER_0_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1620_ _1771_/Q _1620_/B VGND VGND VPWR VPWR _1620_/X sky130_fd_sc_hd__xor2_1
X_1551_ _1708_/A _1818_/Q VGND VGND VPWR VPWR _1551_/Y sky130_fd_sc_hd__nor2_2
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1482_ _1781_/Q _1708_/B VGND VGND VPWR VPWR _1482_/X sky130_fd_sc_hd__or2b_1
XFILLER_39_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1818_ _1818_/D _1668_/C VGND VGND VPWR VPWR _1818_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1749_ _1755_/A _1853_/Q VGND VGND VPWR VPWR _1750_/A sky130_fd_sc_hd__and2_1
XFILLER_53_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0982_ _0999_/A _0997_/A _0997_/B _0974_/X _0980_/A VGND VGND VPWR VPWR _1028_/C
+ sky130_fd_sc_hd__a311o_1
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1603_ _1603_/A _1620_/B VGND VGND VPWR VPWR _1604_/B sky130_fd_sc_hd__xor2_1
X_1534_ _1534_/A _1538_/B VGND VGND VPWR VPWR _1535_/A sky130_fd_sc_hd__and2_1
X_1465_ _1559_/A VGND VGND VPWR VPWR _1523_/A sky130_fd_sc_hd__clkbuf_1
X_1396_ _1396_/A _1396_/B VGND VGND VPWR VPWR _1398_/C sky130_fd_sc_hd__xnor2_1
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1250_ _1388_/A _1347_/A _1249_/B _1335_/A VGND VGND VPWR VPWR _1250_/X sky130_fd_sc_hd__a22o_1
X_1181_ _1181_/A _1212_/A VGND VGND VPWR VPWR _1202_/A sky130_fd_sc_hd__nor2_1
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0965_ _1204_/B _0995_/A _0995_/B VGND VGND VPWR VPWR _0999_/A sky130_fd_sc_hd__or3_1
X_0896_ _1829_/Q VGND VGND VPWR VPWR _0950_/A sky130_fd_sc_hd__clkbuf_1
X_1448_ _1448_/A VGND VGND VPWR VPWR _1448_/Y sky130_fd_sc_hd__inv_2
X_1517_ _1534_/A _1532_/B _1523_/A VGND VGND VPWR VPWR _1518_/A sky130_fd_sc_hd__and3_1
X_1379_ _1447_/B _1379_/B VGND VGND VPWR VPWR _1379_/X sky130_fd_sc_hd__and2_1
XFILLER_23_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1302_ _1334_/B _1302_/B VGND VGND VPWR VPWR _1310_/A sky130_fd_sc_hd__nor2_1
X_1233_ _1263_/A _1233_/B VGND VGND VPWR VPWR _1235_/B sky130_fd_sc_hd__or2_1
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1095_ _0921_/A _1094_/X _1061_/A _1061_/B VGND VGND VPWR VPWR _1146_/B sky130_fd_sc_hd__a211o_1
XFILLER_52_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1164_ input4/X VGND VGND VPWR VPWR _1711_/S sky130_fd_sc_hd__clkbuf_2
X_0948_ _1830_/Q _0983_/B _0983_/C _0947_/Y VGND VGND VPWR VPWR _0968_/C sky130_fd_sc_hd__o31a_2
X_0879_ _1554_/A _1530_/B VGND VGND VPWR VPWR _0880_/A sky130_fd_sc_hd__or2_1
XFILLER_55_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1851_ _1816_/Q _1851_/D VGND VGND VPWR VPWR _1851_/Q sky130_fd_sc_hd__dfxtp_1
X_1782_ _1816_/Q _1782_/D VGND VGND VPWR VPWR _1782_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1216_ _1693_/A VGND VGND VPWR VPWR _1456_/A sky130_fd_sc_hd__buf_2
X_1147_ _1100_/C _1109_/A _1144_/A _1101_/D VGND VGND VPWR VPWR _1147_/Y sky130_fd_sc_hd__a211oi_1
X_1078_ _1133_/A _1070_/A _1070_/B _1123_/A VGND VGND VPWR VPWR _1078_/X sky130_fd_sc_hd__a31o_1
XFILLER_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1001_ _0996_/Y _1000_/Y _1008_/S VGND VGND VPWR VPWR _1024_/B sky130_fd_sc_hd__mux2_1
XFILLER_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1834_ _1834_/D _1666_/A VGND VGND VPWR VPWR _1834_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_30_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1765_ _1816_/Q _1765_/D VGND VGND VPWR VPWR _1765_/Q sky130_fd_sc_hd__dfxtp_1
X_1696_ _1851_/Q _1852_/Q _1696_/C VGND VGND VPWR VPWR _1696_/X sky130_fd_sc_hd__and3_1
XFILLER_13_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput12 _1511_/Y VGND VGND VPWR VPWR seven_segment_out[4] sky130_fd_sc_hd__buf_2
XFILLER_31_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1550_ _1550_/A VGND VGND VPWR VPWR _1826_/D sky130_fd_sc_hd__clkbuf_1
XTAP_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1481_ _1512_/A VGND VGND VPWR VPWR _1485_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_54_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1817_ _1816_/Q _1817_/D VGND VGND VPWR VPWR _1817_/Q sky130_fd_sc_hd__dfxtp_1
X_1748_ _1748_/A VGND VGND VPWR VPWR _1853_/D sky130_fd_sc_hd__clkbuf_1
X_1679_ _1679_/A VGND VGND VPWR VPWR _1688_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_45_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0981_ _0981_/A _0981_/B VGND VGND VPWR VPWR _0981_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_44_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1602_ _1536_/A _1620_/B _1595_/X VGND VGND VPWR VPWR _1604_/A sky130_fd_sc_hd__a21o_1
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1395_ _1347_/Y _1393_/Y _1394_/X VGND VGND VPWR VPWR _1396_/B sky130_fd_sc_hd__o21ai_1
X_1533_ _1533_/A VGND VGND VPWR VPWR _1834_/D sky130_fd_sc_hd__clkbuf_1
X_1464_ _1838_/Q _1665_/A VGND VGND VPWR VPWR _1559_/A sky130_fd_sc_hd__nor2_1
XFILLER_50_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1180_ _1180_/A _1198_/B VGND VGND VPWR VPWR _1212_/A sky130_fd_sc_hd__nand2_1
X_0964_ _1244_/A _1244_/B _0964_/C VGND VGND VPWR VPWR _0995_/B sky130_fd_sc_hd__and3_1
XFILLER_32_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0895_ _1339_/D VGND VGND VPWR VPWR _1388_/C sky130_fd_sc_hd__clkbuf_2
X_1516_ _1516_/A VGND VGND VPWR VPWR _1532_/B sky130_fd_sc_hd__clkbuf_1
X_1378_ _1447_/A _1332_/B _1377_/Y VGND VGND VPWR VPWR _1379_/B sky130_fd_sc_hd__o21ai_1
X_1447_ _1447_/A _1447_/B VGND VGND VPWR VPWR _1447_/Y sky130_fd_sc_hd__nand2_1
XFILLER_11_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1301_ _1299_/C _1341_/B _1300_/Y _1334_/A VGND VGND VPWR VPWR _1302_/B sky130_fd_sc_hd__o2bb2a_1
X_1232_ _1232_/A _1232_/B VGND VGND VPWR VPWR _1233_/B sky130_fd_sc_hd__nor2_1
XFILLER_64_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1094_ _1086_/A _1085_/A _1085_/B _0992_/A VGND VGND VPWR VPWR _1094_/X sky130_fd_sc_hd__a31o_1
XFILLER_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1163_ _1178_/A _1277_/B _1183_/A VGND VGND VPWR VPWR _1163_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_60_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0947_ _0945_/Y _0946_/X _0927_/Y VGND VGND VPWR VPWR _0947_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_20_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0878_ _1516_/A VGND VGND VPWR VPWR _1530_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_28_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1781_ _1816_/Q _1781_/D VGND VGND VPWR VPWR _1781_/Q sky130_fd_sc_hd__dfxtp_1
X_1850_ _1816_/Q _1850_/D VGND VGND VPWR VPWR _1850_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1146_ _1146_/A _1146_/B VGND VGND VPWR VPWR _1146_/Y sky130_fd_sc_hd__nand2_1
XFILLER_25_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1215_ _1727_/B VGND VGND VPWR VPWR _1693_/A sky130_fd_sc_hd__clkbuf_2
X_1077_ _1162_/A _1421_/A VGND VGND VPWR VPWR _1123_/A sky130_fd_sc_hd__nor2_1
XFILLER_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1000_ _1000_/A _1000_/B VGND VGND VPWR VPWR _1000_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1833_ _1833_/D _1666_/A VGND VGND VPWR VPWR _1833_/Q sky130_fd_sc_hd__dlxtn_2
XFILLER_30_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1764_ _1816_/Q _1764_/D VGND VGND VPWR VPWR _1764_/Q sky130_fd_sc_hd__dfxtp_1
X_1695_ _1854_/Q _1855_/Q _1856_/Q _1857_/Q VGND VGND VPWR VPWR _1696_/C sky130_fd_sc_hd__and4_1
X_1129_ _1299_/C VGND VGND VPWR VPWR _1335_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_40_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput13 _1514_/X VGND VGND VPWR VPWR seven_segment_out[5] sky130_fd_sc_hd__buf_2
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1480_ _1498_/B VGND VGND VPWR VPWR _1512_/A sky130_fd_sc_hd__inv_2
XFILLER_47_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1816_ _1839_/CLK _1816_/D VGND VGND VPWR VPWR _1816_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_7_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1747_ _1747_/A _1852_/Q VGND VGND VPWR VPWR _1748_/A sky130_fd_sc_hd__and2_1
X_1678_ _1678_/A VGND VGND VPWR VPWR _1796_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0980_ _0980_/A _1028_/B VGND VGND VPWR VPWR _0981_/B sky130_fd_sc_hd__or2b_1
X_1532_ _1773_/Q _1532_/B _1532_/C VGND VGND VPWR VPWR _1533_/A sky130_fd_sc_hd__and3_1
X_1601_ _1624_/B VGND VGND VPWR VPWR _1620_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_8_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1394_ _1347_/A _1393_/B _1221_/B _1393_/A VGND VGND VPWR VPWR _1394_/X sky130_fd_sc_hd__a22o_1
X_1463_ _1788_/Q _1818_/D _1805_/D _1603_/A VGND VGND VPWR VPWR _1814_/D sky130_fd_sc_hd__a22o_1
XFILLER_35_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0963_ _0968_/A _0963_/B VGND VGND VPWR VPWR _0964_/C sky130_fd_sc_hd__xnor2_1
X_0894_ _0985_/A VGND VGND VPWR VPWR _1339_/D sky130_fd_sc_hd__clkbuf_2
X_1515_ _1491_/X _1485_/A _1505_/B _1499_/B VGND VGND VPWR VPWR _1515_/X sky130_fd_sc_hd__a211o_1
X_1446_ _1446_/A _1446_/B VGND VGND VPWR VPWR _1446_/Y sky130_fd_sc_hd__nand2_1
X_1377_ _1420_/A _1422_/B VGND VGND VPWR VPWR _1377_/Y sky130_fd_sc_hd__nand2_1
XFILLER_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1300_ _1300_/A VGND VGND VPWR VPWR _1300_/Y sky130_fd_sc_hd__clkinv_2
X_1162_ _1162_/A _1382_/A VGND VGND VPWR VPWR _1277_/B sky130_fd_sc_hd__and2_1
XFILLER_37_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1231_ _1232_/A _1232_/B VGND VGND VPWR VPWR _1263_/A sky130_fd_sc_hd__and2_1
XFILLER_1_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1093_ _1093_/A VGND VGND VPWR VPWR _1146_/A sky130_fd_sc_hd__inv_2
XFILLER_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0946_ _0956_/A _0946_/B _0946_/C VGND VGND VPWR VPWR _0946_/X sky130_fd_sc_hd__and3_1
X_0877_ _1837_/Q VGND VGND VPWR VPWR _1516_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1429_ _1376_/A _1137_/A _1426_/X _1427_/Y VGND VGND VPWR VPWR _1429_/X sky130_fd_sc_hd__a211o_1
XFILLER_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1780_ _1816_/Q _1780_/D VGND VGND VPWR VPWR _1780_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1145_ _1141_/X _1144_/Y _1149_/S VGND VGND VPWR VPWR _1145_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1214_ _1212_/X _1222_/A _1193_/X VGND VGND VPWR VPWR _1214_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_25_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1076_ _1180_/A VGND VGND VPWR VPWR _1421_/A sky130_fd_sc_hd__clkbuf_2
X_0929_ _0945_/A _0945_/B _0935_/C VGND VGND VPWR VPWR _1287_/A sky130_fd_sc_hd__and3_1
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1832_ _1832_/D _1666_/A VGND VGND VPWR VPWR _1832_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_42_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1694_ _1694_/A VGND VGND VPWR VPWR _1851_/D sky130_fd_sc_hd__clkbuf_1
X_1763_ _1816_/Q _1763_/D VGND VGND VPWR VPWR _1763_/Q sky130_fd_sc_hd__dfxtp_1
X_1059_ _1022_/X _1059_/B VGND VGND VPWR VPWR _1060_/B sky130_fd_sc_hd__and2b_1
X_1128_ _1819_/Q VGND VGND VPWR VPWR _1299_/C sky130_fd_sc_hd__clkbuf_1
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput14 _1515_/X VGND VGND VPWR VPWR seven_segment_out[6] sky130_fd_sc_hd__buf_2
XFILLER_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1815_ _1815_/D _1667_/B VGND VGND VPWR VPWR _1815_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_7_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1746_ _1746_/A VGND VGND VPWR VPWR _1852_/D sky130_fd_sc_hd__clkbuf_1
X_1677_ _1693_/A _1795_/Q VGND VGND VPWR VPWR _1678_/A sky130_fd_sc_hd__and2_1
XFILLER_26_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1531_ _1531_/A VGND VGND VPWR VPWR _1833_/D sky130_fd_sc_hd__clkbuf_1
X_1600_ _1536_/A _1588_/X _1597_/Y _1599_/X VGND VGND VPWR VPWR _1767_/D sky130_fd_sc_hd__o211a_1
X_1462_ _1768_/Q VGND VGND VPWR VPWR _1603_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_8_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1393_ _1393_/A _1393_/B VGND VGND VPWR VPWR _1393_/Y sky130_fd_sc_hd__nand2_1
XFILLER_35_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1729_ _1844_/Q _1735_/B VGND VGND VPWR VPWR _1730_/A sky130_fd_sc_hd__and2_1
XFILLER_58_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0962_ _0961_/X _0962_/B VGND VGND VPWR VPWR _0963_/B sky130_fd_sc_hd__and2b_1
X_0893_ _1831_/Q VGND VGND VPWR VPWR _0985_/A sky130_fd_sc_hd__buf_2
X_1445_ _1445_/A _1445_/B VGND VGND VPWR VPWR _1445_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1514_ _1485_/A _1493_/X _1500_/Y _1513_/X VGND VGND VPWR VPWR _1514_/X sky130_fd_sc_hd__a31o_4
XFILLER_55_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1376_ _1376_/A _1376_/B VGND VGND VPWR VPWR _1447_/B sky130_fd_sc_hd__xnor2_2
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1092_ _1335_/B VGND VGND VPWR VPWR _1411_/B sky130_fd_sc_hd__inv_2
X_1230_ _1257_/B _1230_/B VGND VGND VPWR VPWR _1232_/B sky130_fd_sc_hd__nor2_1
XFILLER_37_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1161_ _1154_/X _1157_/Y _1315_/A _1179_/B _1183_/A VGND VGND VPWR VPWR _1161_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_1_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0945_ _0945_/A _0945_/B VGND VGND VPWR VPWR _0945_/Y sky130_fd_sc_hd__nand2_1
X_0876_ _1668_/B VGND VGND VPWR VPWR _1554_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_9_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1428_ _1426_/X _1427_/Y _1137_/A VGND VGND VPWR VPWR _1428_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1359_ _1360_/A _1360_/B _1360_/C VGND VGND VPWR VPWR _1381_/A sky130_fd_sc_hd__a21oi_1
XFILLER_28_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1213_ _1212_/A _1212_/B _1207_/A VGND VGND VPWR VPWR _1222_/A sky130_fd_sc_hd__a21oi_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1144_ _1144_/A _1144_/B VGND VGND VPWR VPWR _1144_/Y sky130_fd_sc_hd__xnor2_1
X_1075_ _1341_/C VGND VGND VPWR VPWR _1180_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_37_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0928_ _0956_/A _0946_/B _0946_/C _0927_/Y VGND VGND VPWR VPWR _0935_/C sky130_fd_sc_hd__a31o_1
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1831_ _1831_/D _1666_/A VGND VGND VPWR VPWR _1831_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_15_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1693_ _1693_/A _1850_/Q VGND VGND VPWR VPWR _1694_/A sky130_fd_sc_hd__and2_1
X_1762_ _1816_/Q _1762_/D VGND VGND VPWR VPWR _1762_/Q sky130_fd_sc_hd__dfxtp_1
X_1058_ _1058_/A VGND VGND VPWR VPWR _1058_/Y sky130_fd_sc_hd__inv_2
X_1127_ _1820_/Q VGND VGND VPWR VPWR _1197_/A sky130_fd_sc_hd__inv_2
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1745_ _1747_/A _1851_/Q VGND VGND VPWR VPWR _1746_/A sky130_fd_sc_hd__and2_1
X_1814_ _1814_/D _1667_/B VGND VGND VPWR VPWR _1814_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1676_ _1676_/A VGND VGND VPWR VPWR _1795_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_53_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1392_ _1392_/A _1392_/B VGND VGND VPWR VPWR _1396_/A sky130_fd_sc_hd__nor2_1
X_1530_ _1547_/A _1530_/B _1532_/C VGND VGND VPWR VPWR _1531_/A sky130_fd_sc_hd__and3_1
X_1461_ _1787_/Q _1818_/D _1805_/D _1536_/A VGND VGND VPWR VPWR _1813_/D sky130_fd_sc_hd__a22o_1
XFILLER_50_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1728_ _1728_/A VGND VGND VPWR VPWR _1844_/D sky130_fd_sc_hd__clkbuf_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1659_ _1781_/Q _1811_/Q _1805_/Q VGND VGND VPWR VPWR _1660_/B sky130_fd_sc_hd__mux2_1
XFILLER_41_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0961_ _1350_/B _0961_/B _0961_/C VGND VGND VPWR VPWR _0961_/X sky130_fd_sc_hd__and3_1
XFILLER_17_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0892_ _1426_/B VGND VGND VPWR VPWR _1290_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_40_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1375_ _1826_/Q VGND VGND VPWR VPWR _1376_/A sky130_fd_sc_hd__buf_2
X_1444_ _1444_/A _1444_/B VGND VGND VPWR VPWR _1445_/B sky130_fd_sc_hd__xnor2_1
X_1513_ _1491_/X _1505_/A _1505_/B _1499_/B _1512_/X VGND VGND VPWR VPWR _1513_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1091_ _1833_/Q VGND VGND VPWR VPWR _1335_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_45_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1160_ _1807_/Q VGND VGND VPWR VPWR _1183_/A sky130_fd_sc_hd__inv_2
X_0944_ _0950_/A _0951_/B _0962_/B _0949_/B VGND VGND VPWR VPWR _0983_/C sky130_fd_sc_hd__o211a_1
XFILLER_9_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0875_ _1838_/Q VGND VGND VPWR VPWR _1668_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1358_ _1402_/B _1358_/B VGND VGND VPWR VPWR _1360_/C sky130_fd_sc_hd__nand2_1
X_1427_ _1426_/A _1290_/B _1426_/C VGND VGND VPWR VPWR _1427_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1289_ _1289_/A VGND VGND VPWR VPWR _1291_/A sky130_fd_sc_hd__inv_2
XFILLER_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1212_ _1212_/A _1212_/B _1276_/A VGND VGND VPWR VPWR _1212_/X sky130_fd_sc_hd__and3_1
X_1143_ _1100_/C _1109_/A _1101_/D VGND VGND VPWR VPWR _1144_/B sky130_fd_sc_hd__a21o_1
X_1074_ _1820_/Q VGND VGND VPWR VPWR _1341_/C sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0927_ _0937_/A _0926_/Y _0902_/X VGND VGND VPWR VPWR _0927_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1830_ _1830_/D _1666_/A VGND VGND VPWR VPWR _1830_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_15_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1761_ _1816_/Q _1761_/D VGND VGND VPWR VPWR _1761_/Q sky130_fd_sc_hd__dfxtp_1
X_1692_ _1692_/A VGND VGND VPWR VPWR _1802_/D sky130_fd_sc_hd__clkbuf_1
X_1126_ _1420_/B _1126_/B _1126_/C VGND VGND VPWR VPWR _1126_/X sky130_fd_sc_hd__or3_1
X_1057_ _1057_/A _1057_/B VGND VGND VPWR VPWR _1058_/A sky130_fd_sc_hd__and2_1
XFILLER_40_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1813_ _1813_/D _1667_/B VGND VGND VPWR VPWR _1813_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1744_ _1744_/A VGND VGND VPWR VPWR _1850_/D sky130_fd_sc_hd__clkbuf_1
X_1675_ _1675_/A input2/X VGND VGND VPWR VPWR _1676_/A sky130_fd_sc_hd__and2_1
X_1109_ _1109_/A _1109_/B VGND VGND VPWR VPWR _1109_/Y sky130_fd_sc_hd__nand2_1
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1391_ _1391_/A _1391_/B VGND VGND VPWR VPWR _1400_/A sky130_fd_sc_hd__xor2_2
X_1460_ _1807_/D VGND VGND VPWR VPWR _1536_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_50_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1727_ _1843_/Q _1727_/B VGND VGND VPWR VPWR _1728_/A sky130_fd_sc_hd__and2_1
X_1658_ _1658_/A VGND VGND VPWR VPWR _1780_/D sky130_fd_sc_hd__clkbuf_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1589_ _1534_/A _1596_/A _1711_/S VGND VGND VPWR VPWR _1589_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_53_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0960_ _1348_/C _0983_/B _0983_/C _0947_/Y VGND VGND VPWR VPWR _1244_/B sky130_fd_sc_hd__o31ai_2
XFILLER_32_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0891_ _1387_/B VGND VGND VPWR VPWR _1426_/B sky130_fd_sc_hd__clkbuf_2
X_1512_ _1512_/A _1512_/B _1512_/C VGND VGND VPWR VPWR _1512_/X sky130_fd_sc_hd__and3_1
XFILLER_55_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1443_ _1443_/A _1443_/B VGND VGND VPWR VPWR _1444_/B sky130_fd_sc_hd__xnor2_1
X_1374_ _1193_/X _1332_/Y _1373_/X _1708_/A VGND VGND VPWR VPWR _1792_/D sky130_fd_sc_hd__a211oi_1
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1090_ _1061_/A _1061_/B _1086_/X _1089_/X _1387_/B VGND VGND VPWR VPWR _1142_/B
+ sky130_fd_sc_hd__o311a_1
XFILLER_38_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0943_ _0950_/A _0951_/B VGND VGND VPWR VPWR _0983_/B sky130_fd_sc_hd__and2_1
XFILLER_9_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1357_ _1357_/A _1357_/B VGND VGND VPWR VPWR _1358_/B sky130_fd_sc_hd__or2_1
X_1426_ _1426_/A _1426_/B _1426_/C VGND VGND VPWR VPWR _1426_/X sky130_fd_sc_hd__and3_1
X_1288_ _1290_/A _1426_/B VGND VGND VPWR VPWR _1289_/A sky130_fd_sc_hd__nand2_1
XFILLER_28_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1142_ _1142_/A _1142_/B VGND VGND VPWR VPWR _1144_/A sky130_fd_sc_hd__or2_1
X_1211_ _1195_/X _1245_/A _1203_/X _1209_/X _1210_/X VGND VGND VPWR VPWR _1211_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1073_ _1198_/B VGND VGND VPWR VPWR _1133_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_33_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0926_ _0902_/X _0904_/X _0907_/X VGND VGND VPWR VPWR _0926_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1409_ _1409_/A _1409_/B _1409_/C VGND VGND VPWR VPWR _1409_/X sky130_fd_sc_hd__or3_1
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1691_ _1747_/A _1801_/Q VGND VGND VPWR VPWR _1692_/A sky130_fd_sc_hd__and2_1
X_1760_ _1816_/Q _1760_/D VGND VGND VPWR VPWR _1760_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1125_ _1114_/B _1124_/S _1119_/X _1220_/B VGND VGND VPWR VPWR _1126_/C sky130_fd_sc_hd__o211a_1
XFILLER_25_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1056_ _1107_/A _1107_/B _1112_/A VGND VGND VPWR VPWR _1101_/A sky130_fd_sc_hd__a21oi_1
XFILLER_40_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0909_ _0902_/X _0904_/X _0907_/X _0966_/A VGND VGND VPWR VPWR _0910_/B sky130_fd_sc_hd__a211o_1
XFILLER_31_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1674_ _1785_/Q _1668_/X _1672_/X _1673_/Y VGND VGND VPWR VPWR _1785_/D sky130_fd_sc_hd__a22o_1
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1743_ _1747_/A input3/X VGND VGND VPWR VPWR _1744_/A sky130_fd_sc_hd__and2_1
X_1812_ _1812_/D _1667_/B VGND VGND VPWR VPWR _1812_/Q sky130_fd_sc_hd__dlxtn_1
X_1108_ _1116_/A _1082_/B _1082_/C VGND VGND VPWR VPWR _1109_/B sky130_fd_sc_hd__o21ai_1
X_1039_ _1039_/A VGND VGND VPWR VPWR _1085_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1390_ _1826_/Q _1388_/X _1389_/X VGND VGND VPWR VPWR _1391_/B sky130_fd_sc_hd__a21bo_1
XFILLER_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1588_ _1596_/A VGND VGND VPWR VPWR _1588_/X sky130_fd_sc_hd__clkbuf_2
X_1726_ _1726_/A VGND VGND VPWR VPWR _1843_/D sky130_fd_sc_hd__clkbuf_1
X_1657_ _1675_/A _1657_/B VGND VGND VPWR VPWR _1658_/A sky130_fd_sc_hd__and2_1
XFILLER_58_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0890_ _1341_/B VGND VGND VPWR VPWR _1387_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_43_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1442_ _1442_/A _1442_/B VGND VGND VPWR VPWR _1443_/B sky130_fd_sc_hd__xnor2_1
X_1511_ _1511_/A _1511_/B VGND VGND VPWR VPWR _1511_/Y sky130_fd_sc_hd__nand2_4
X_1373_ _1409_/B _1369_/X _1372_/Y VGND VGND VPWR VPWR _1373_/X sky130_fd_sc_hd__o21a_1
XFILLER_4_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1709_ _1783_/Q _1665_/A _1711_/S VGND VGND VPWR VPWR _1710_/A sky130_fd_sc_hd__mux2_1
XFILLER_64_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0942_ _1830_/Q _0932_/X _0941_/X _0985_/A _0907_/B VGND VGND VPWR VPWR _0968_/B
+ sky130_fd_sc_hd__a311o_2
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1425_ _1425_/A _1425_/B VGND VGND VPWR VPWR _1431_/A sky130_fd_sc_hd__xnor2_1
XFILLER_55_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1356_ _1357_/A _1357_/B VGND VGND VPWR VPWR _1402_/B sky130_fd_sc_hd__nand2_1
X_1287_ _1287_/A _1287_/B VGND VGND VPWR VPWR _1287_/X sky130_fd_sc_hd__and2_1
XFILLER_36_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1141_ _1062_/S _1086_/X _1087_/X VGND VGND VPWR VPWR _1141_/X sky130_fd_sc_hd__a21o_1
X_1072_ _1304_/B VGND VGND VPWR VPWR _1198_/B sky130_fd_sc_hd__clkbuf_2
X_1210_ _1210_/A VGND VGND VPWR VPWR _1210_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0925_ _0946_/B _0946_/C _0956_/A VGND VGND VPWR VPWR _0945_/B sky130_fd_sc_hd__a21o_1
X_1408_ _1408_/A _1408_/B VGND VGND VPWR VPWR _1409_/C sky130_fd_sc_hd__xor2_1
XFILLER_29_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1339_ _1339_/A _1420_/A _1387_/A _1339_/D VGND VGND VPWR VPWR _1339_/X sky130_fd_sc_hd__and4_1
XFILLER_45_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1690_ _1690_/A VGND VGND VPWR VPWR _1747_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1055_ _1055_/A _1069_/A _1069_/C _1055_/D VGND VGND VPWR VPWR _1107_/B sky130_fd_sc_hd__or4_1
X_1124_ _1122_/B _1123_/Y _1124_/S VGND VGND VPWR VPWR _1126_/B sky130_fd_sc_hd__mux2_1
XFILLER_53_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0908_ _1827_/Q VGND VGND VPWR VPWR _0966_/A sky130_fd_sc_hd__inv_2
XFILLER_0_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1811_ _1811_/D _1667_/B VGND VGND VPWR VPWR _1811_/Q sky130_fd_sc_hd__dlxtn_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1673_ _1849_/Q VGND VGND VPWR VPWR _1673_/Y sky130_fd_sc_hd__inv_2
XFILLER_7_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1742_ _1737_/X _1738_/X _1741_/X VGND VGND VPWR VPWR _1849_/D sky130_fd_sc_hd__o21a_1
X_1107_ _1107_/A _1107_/B VGND VGND VPWR VPWR _1107_/X sky130_fd_sc_hd__and2_1
X_1038_ _1061_/A _1061_/B _1024_/B VGND VGND VPWR VPWR _1047_/B sky130_fd_sc_hd__o21ai_1
XFILLER_53_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1725_ _1842_/Q _1725_/B VGND VGND VPWR VPWR _1726_/A sky130_fd_sc_hd__and2_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1587_ _1609_/C VGND VGND VPWR VPWR _1596_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1656_ _1780_/Q _1810_/Q _1805_/Q VGND VGND VPWR VPWR _1657_/B sky130_fd_sc_hd__mux2_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1441_ _1396_/A _1394_/X _1393_/Y _1440_/Y VGND VGND VPWR VPWR _1442_/B sky130_fd_sc_hd__a31o_1
XFILLER_4_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1510_ _1493_/X _1504_/A _1491_/X VGND VGND VPWR VPWR _1511_/B sky130_fd_sc_hd__a21bo_1
XFILLER_48_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1372_ _0926_/Y _1171_/A _1210_/X _1371_/Y _1193_/A VGND VGND VPWR VPWR _1372_/Y
+ sky130_fd_sc_hd__a221oi_2
XFILLER_63_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1708_ _1708_/A _1708_/B VGND VGND VPWR VPWR _1835_/D sky130_fd_sc_hd__nor2_1
XFILLER_2_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1639_ _1639_/A VGND VGND VPWR VPWR _1774_/D sky130_fd_sc_hd__clkbuf_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0941_ _0950_/A _0931_/A _0962_/B _0949_/B VGND VGND VPWR VPWR _0941_/X sky130_fd_sc_hd__a22o_1
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1424_ _1424_/A _1424_/B VGND VGND VPWR VPWR _1425_/B sky130_fd_sc_hd__xnor2_1
X_1355_ _1402_/A _1355_/B VGND VGND VPWR VPWR _1357_/B sky130_fd_sc_hd__and2_1
XFILLER_55_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1286_ _1193_/X _1244_/X _1280_/X _1285_/X _1217_/X VGND VGND VPWR VPWR _1790_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_63_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1071_ _1350_/B VGND VGND VPWR VPWR _1304_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_45_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1140_ _1335_/B VGND VGND VPWR VPWR _1422_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_37_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0924_ _1829_/Q VGND VGND VPWR VPWR _0956_/A sky130_fd_sc_hd__inv_2
XFILLER_33_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1407_ _1407_/A _1437_/A VGND VGND VPWR VPWR _1408_/B sky130_fd_sc_hd__xor2_1
X_1338_ _1338_/A _1308_/B VGND VGND VPWR VPWR _1360_/A sky130_fd_sc_hd__or2b_1
XFILLER_45_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1269_ _1270_/A _1270_/B VGND VGND VPWR VPWR _1271_/A sky130_fd_sc_hd__nor2_1
XFILLER_24_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1054_ _1054_/A _1054_/B VGND VGND VPWR VPWR _1055_/D sky130_fd_sc_hd__and2_1
X_1123_ _1123_/A _1123_/B VGND VGND VPWR VPWR _1123_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_25_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0907_ _1829_/Q _0907_/B _0907_/C _0921_/B VGND VGND VPWR VPWR _0907_/X sky130_fd_sc_hd__or4b_1
XFILLER_56_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1810_ _1810_/D _1667_/B VGND VGND VPWR VPWR _1810_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1741_ _1844_/D _1739_/X _1740_/X _1456_/A _1849_/Q VGND VGND VPWR VPWR _1741_/X
+ sky130_fd_sc_hd__a32o_1
X_1672_ _0883_/A _0887_/X _1672_/S VGND VGND VPWR VPWR _1672_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1106_ _1044_/Y _1084_/Y _1149_/S VGND VGND VPWR VPWR _1106_/X sky130_fd_sc_hd__mux2_1
X_1037_ _1069_/C VGND VGND VPWR VPWR _1061_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1724_ _1724_/A VGND VGND VPWR VPWR _1842_/D sky130_fd_sc_hd__clkbuf_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1586_ _1582_/X _1583_/X _1584_/X _1585_/Y VGND VGND VPWR VPWR _1609_/C sky130_fd_sc_hd__o22a_1
X_1655_ _1655_/A VGND VGND VPWR VPWR _1779_/D sky130_fd_sc_hd__clkbuf_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1440_ _1270_/A _1420_/B _1396_/A _1394_/X _1393_/Y VGND VGND VPWR VPWR _1440_/Y
+ sky130_fd_sc_hd__a221oi_1
X_1371_ _1447_/A _1371_/B VGND VGND VPWR VPWR _1371_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1638_ _1647_/A _1638_/B VGND VGND VPWR VPWR _1639_/A sky130_fd_sc_hd__and2_1
X_1707_ _1797_/Q _1796_/D _1703_/X _1706_/X VGND VGND VPWR VPWR _1817_/D sky130_fd_sc_hd__a31o_1
XFILLER_39_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1569_ _1759_/Q _1693_/A VGND VGND VPWR VPWR _1570_/A sky130_fd_sc_hd__and2_1
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0940_ _0937_/A _0961_/B _0961_/C _0968_/A VGND VGND VPWR VPWR _0949_/B sky130_fd_sc_hd__a31o_1
X_1423_ _1423_/A _1423_/B VGND VGND VPWR VPWR _1424_/B sky130_fd_sc_hd__xor2_1
X_1354_ _1354_/A _1354_/B _1354_/C VGND VGND VPWR VPWR _1355_/B sky130_fd_sc_hd__or3_1
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1285_ _1283_/Y _1323_/B _1193_/A VGND VGND VPWR VPWR _1285_/X sky130_fd_sc_hd__a21bo_1
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1070_ _1070_/A _1070_/B VGND VGND VPWR VPWR _1122_/B sky130_fd_sc_hd__and2_1
XFILLER_52_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0923_ _1327_/A _1020_/A _0910_/B _1350_/A _0966_/A VGND VGND VPWR VPWR _0946_/C
+ sky130_fd_sc_hd__a311o_1
XFILLER_33_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1337_ _1407_/A _1337_/B VGND VGND VPWR VPWR _1361_/A sky130_fd_sc_hd__or2_1
X_1406_ _1438_/A _1438_/B VGND VGND VPWR VPWR _1437_/A sky130_fd_sc_hd__xnor2_1
X_1268_ _1268_/A _1268_/B VGND VGND VPWR VPWR _1268_/Y sky130_fd_sc_hd__nand2_1
XFILLER_28_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1199_ _1212_/A _1225_/A _1232_/A VGND VGND VPWR VPWR _1201_/B sky130_fd_sc_hd__a21o_1
XFILLER_24_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1122_ _1133_/A _1122_/B VGND VGND VPWR VPWR _1123_/B sky130_fd_sc_hd__xnor2_1
X_1053_ _1054_/A _1054_/B VGND VGND VPWR VPWR _1055_/A sky130_fd_sc_hd__nor2_1
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0906_ _1825_/Q _1828_/Q _1827_/Q VGND VGND VPWR VPWR _0907_/C sky130_fd_sc_hd__and3b_1
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1671_ _1784_/Q _1668_/X _1670_/X _1667_/Y VGND VGND VPWR VPWR _1784_/D sky130_fd_sc_hd__a22o_1
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1740_ _1842_/Q _1841_/Q _1844_/Q _1846_/Q VGND VGND VPWR VPWR _1740_/X sky130_fd_sc_hd__and4_1
XFILLER_15_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1105_ _1124_/S VGND VGND VPWR VPWR _1149_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_38_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1036_ _1051_/A _1051_/B VGND VGND VPWR VPWR _1069_/C sky130_fd_sc_hd__nand2_1
XFILLER_29_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1723_ _1841_/Q _1725_/B VGND VGND VPWR VPWR _1724_/A sky130_fd_sc_hd__and2_1
X_1654_ _1675_/A _1654_/B VGND VGND VPWR VPWR _1655_/A sky130_fd_sc_hd__and2_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1585_ _1782_/Q _1757_/Q VGND VGND VPWR VPWR _1585_/Y sky130_fd_sc_hd__nor2_1
X_1019_ _1235_/A _1018_/X _0988_/A _0988_/B VGND VGND VPWR VPWR _1057_/B sky130_fd_sc_hd__a211o_1
XFILLER_34_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1370_ _1289_/A _1294_/B _1291_/B VGND VGND VPWR VPWR _1371_/B sky130_fd_sc_hd__a21oi_1
XFILLER_23_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1637_ _1774_/Q _1812_/Q _1650_/S VGND VGND VPWR VPWR _1638_/B sky130_fd_sc_hd__mux2_1
X_1706_ _1704_/X _1705_/X _1817_/Q _1456_/A VGND VGND VPWR VPWR _1706_/X sky130_fd_sc_hd__o211a_1
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1499_ _1500_/A _1499_/B VGND VGND VPWR VPWR _1507_/A sky130_fd_sc_hd__and2_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1568_ _1568_/A VGND VGND VPWR VPWR _1759_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_54_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1422_ _1422_/A _1422_/B VGND VGND VPWR VPWR _1423_/B sky130_fd_sc_hd__nand2_1
X_1353_ _1354_/A _1354_/B _1354_/C VGND VGND VPWR VPWR _1402_/A sky130_fd_sc_hd__o21ai_1
X_1284_ _1283_/A _1345_/B _1446_/A VGND VGND VPWR VPWR _1323_/B sky130_fd_sc_hd__a21o_1
XFILLER_51_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0999_ _0999_/A _0999_/B VGND VGND VPWR VPWR _1000_/B sky130_fd_sc_hd__nand2_1
XFILLER_59_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0922_ _1824_/Q VGND VGND VPWR VPWR _1350_/A sky130_fd_sc_hd__clkbuf_2
X_1405_ _1405_/A _1405_/B VGND VGND VPWR VPWR _1438_/B sky130_fd_sc_hd__nor2_1
X_1336_ _1335_/A _1335_/B _1335_/C VGND VGND VPWR VPWR _1337_/B sky130_fd_sc_hd__a21oi_1
X_1198_ _1299_/C _1198_/B _1253_/C VGND VGND VPWR VPWR _1232_/A sky130_fd_sc_hd__and3_1
X_1267_ _1268_/A _1268_/B VGND VGND VPWR VPWR _1320_/A sky130_fd_sc_hd__or2_1
Xinput1 restart VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_36_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1052_ _1194_/A _1194_/B _1026_/B VGND VGND VPWR VPWR _1107_/A sky130_fd_sc_hd__a21o_1
X_1121_ _1220_/B _1121_/B VGND VGND VPWR VPWR _1121_/X sky130_fd_sc_hd__or2_1
XFILLER_33_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0905_ _1833_/Q _1832_/Q _1834_/Q VGND VGND VPWR VPWR _0907_/B sky130_fd_sc_hd__or3_2
XFILLER_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1319_ _1319_/A _1319_/B VGND VGND VPWR VPWR _1320_/B sky130_fd_sc_hd__xor2_1
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1670_ _1538_/B _1672_/S _1666_/Y _1516_/A VGND VGND VPWR VPWR _1670_/X sky130_fd_sc_hd__a22o_1
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1104_ _1100_/X _1103_/X _1421_/B VGND VGND VPWR VPWR _1124_/S sky130_fd_sc_hd__a21oi_2
X_1035_ _1387_/B _1093_/A VGND VGND VPWR VPWR _1051_/B sky130_fd_sc_hd__nand2_1
XFILLER_46_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1799_ _1816_/Q _1799_/D VGND VGND VPWR VPWR _1799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1584_ _1782_/Q _1757_/Q VGND VGND VPWR VPWR _1584_/X sky130_fd_sc_hd__and2_1
XFILLER_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1722_ _1722_/A VGND VGND VPWR VPWR _1841_/D sky130_fd_sc_hd__clkbuf_1
X_1653_ _1779_/Q _1809_/Q _1805_/Q VGND VGND VPWR VPWR _1654_/B sky130_fd_sc_hd__mux2_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1018_ _1018_/A _1822_/Q VGND VGND VPWR VPWR _1018_/X sky130_fd_sc_hd__or2_1
XFILLER_34_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1705_ _1800_/Q _1799_/Q _1801_/Q _1802_/Q VGND VGND VPWR VPWR _1705_/X sky130_fd_sc_hd__or4_1
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1567_ _1758_/Q _1575_/B VGND VGND VPWR VPWR _1568_/A sky130_fd_sc_hd__and2_1
X_1636_ _1805_/Q VGND VGND VPWR VPWR _1650_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_54_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1498_ _1494_/X _1498_/B _1498_/C VGND VGND VPWR VPWR _1499_/B sky130_fd_sc_hd__and3b_1
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1421_ _1421_/A _1421_/B VGND VGND VPWR VPWR _1423_/A sky130_fd_sc_hd__nand2_1
X_1352_ _1398_/B _1352_/B VGND VGND VPWR VPWR _1354_/C sky130_fd_sc_hd__nor2_1
X_1283_ _1283_/A _1446_/A _1345_/B VGND VGND VPWR VPWR _1283_/Y sky130_fd_sc_hd__nand3_1
XFILLER_36_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0998_ _1204_/B _0998_/B VGND VGND VPWR VPWR _0999_/B sky130_fd_sc_hd__nand2_1
XFILLER_59_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1619_ _1614_/A _1616_/B _1613_/Y VGND VGND VPWR VPWR _1619_/X sky130_fd_sc_hd__o21a_1
XFILLER_54_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0921_ _0921_/A _0921_/B VGND VGND VPWR VPWR _0945_/A sky130_fd_sc_hd__and2_1
XFILLER_18_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1404_ _1403_/B _1403_/C _1403_/A VGND VGND VPWR VPWR _1405_/B sky130_fd_sc_hd__a21oi_1
X_1335_ _1335_/A _1335_/B _1335_/C VGND VGND VPWR VPWR _1407_/A sky130_fd_sc_hd__and3_1
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput2 rotary_a VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__clkbuf_2
XFILLER_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1197_ _1197_/A _1204_/B VGND VGND VPWR VPWR _1253_/C sky130_fd_sc_hd__nor2_1
XFILLER_36_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1266_ _1318_/B _1266_/B VGND VGND VPWR VPWR _1268_/B sky130_fd_sc_hd__nand2_1
XFILLER_19_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1120_ _1114_/B _1124_/S _1119_/X VGND VGND VPWR VPWR _1121_/B sky130_fd_sc_hd__o21a_1
X_1051_ _1051_/A _1051_/B VGND VGND VPWR VPWR _1194_/B sky130_fd_sc_hd__and2_1
X_0904_ _1827_/Q _1392_/A _1828_/Q VGND VGND VPWR VPWR _0904_/X sky130_fd_sc_hd__a21o_1
XFILLER_33_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1318_ _1318_/A _1318_/B VGND VGND VPWR VPWR _1319_/B sky130_fd_sc_hd__nand2_1
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1249_ _1270_/A _1249_/B VGND VGND VPWR VPWR _1295_/A sky130_fd_sc_hd__nand2_1
XFILLER_24_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1103_ _1116_/A _1082_/B _1100_/A _1101_/X _1102_/Y VGND VGND VPWR VPWR _1103_/X
+ sky130_fd_sc_hd__o41a_1
X_1034_ _1833_/Q _1421_/B VGND VGND VPWR VPWR _1051_/A sky130_fd_sc_hd__nor2_1
XFILLER_38_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1798_ _1816_/Q _1798_/D VGND VGND VPWR VPWR _1798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1721_ _1747_/A input1/X VGND VGND VPWR VPWR _1722_/A sky130_fd_sc_hd__and2_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1652_ _1652_/A VGND VGND VPWR VPWR _1778_/D sky130_fd_sc_hd__clkbuf_1
X_1583_ _1803_/Q _1817_/Q VGND VGND VPWR VPWR _1583_/X sky130_fd_sc_hd__and2b_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1017_ _1018_/A _1388_/B VGND VGND VPWR VPWR _1235_/A sky130_fd_sc_hd__nand2_2
XFILLER_26_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1704_ _1796_/Q _1795_/Q _1797_/Q _1798_/Q VGND VGND VPWR VPWR _1704_/X sky130_fd_sc_hd__or4_1
XFILLER_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1635_ _1635_/A VGND VGND VPWR VPWR _1773_/D sky130_fd_sc_hd__clkbuf_1
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1497_ _1485_/Y _1492_/X _1496_/Y _1485_/A VGND VGND VPWR VPWR _1497_/X sky130_fd_sc_hd__a22o_2
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1566_ _1566_/A VGND VGND VPWR VPWR _1758_/D sky130_fd_sc_hd__clkbuf_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1420_ _1420_/A _1420_/B VGND VGND VPWR VPWR _1424_/A sky130_fd_sc_hd__nand2_1
X_1351_ _1350_/A _1304_/B _1350_/C VGND VGND VPWR VPWR _1352_/B sky130_fd_sc_hd__a21oi_1
XFILLER_51_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1282_ _1822_/Q _1282_/B VGND VGND VPWR VPWR _1345_/B sky130_fd_sc_hd__nand2_2
XFILLER_36_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0997_ _0997_/A _0997_/B VGND VGND VPWR VPWR _1000_/A sky130_fd_sc_hd__nand2_1
X_1618_ _1613_/A _1588_/X _1617_/Y _1599_/X VGND VGND VPWR VPWR _1770_/D sky130_fd_sc_hd__o211a_1
XFILLER_46_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1549_ _1773_/Q _1549_/B VGND VGND VPWR VPWR _1550_/A sky130_fd_sc_hd__and2_1
XFILLER_54_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0920_ _0920_/A _0920_/B VGND VGND VPWR VPWR _0920_/X sky130_fd_sc_hd__or2_1
XFILLER_45_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1403_ _1403_/A _1403_/B _1403_/C VGND VGND VPWR VPWR _1405_/A sky130_fd_sc_hd__and3_1
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1334_ _1334_/A _1334_/B VGND VGND VPWR VPWR _1335_/C sky130_fd_sc_hd__or2_1
X_1265_ _1318_/A _1264_/C _1246_/X VGND VGND VPWR VPWR _1266_/B sky130_fd_sc_hd__a21bo_1
XFILLER_5_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1196_ _1299_/C _1221_/B VGND VGND VPWR VPWR _1225_/A sky130_fd_sc_hd__nand2_1
Xinput3 rotary_b VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__clkbuf_1
XFILLER_59_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1050_ _1086_/A _1085_/A _1085_/B _0992_/A _1030_/Y VGND VGND VPWR VPWR _1194_/A
+ sky130_fd_sc_hd__a311o_1
XFILLER_33_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0903_ _1825_/Q VGND VGND VPWR VPWR _1392_/A sky130_fd_sc_hd__clkinv_2
XFILLER_33_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1248_ _1347_/A VGND VGND VPWR VPWR _1270_/A sky130_fd_sc_hd__clkbuf_2
X_1317_ _1317_/A _1317_/B VGND VGND VPWR VPWR _1319_/A sky130_fd_sc_hd__or2_1
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1179_ _1807_/Q _1179_/B VGND VGND VPWR VPWR _1210_/A sky130_fd_sc_hd__nor2_1
XFILLER_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1102_ _1142_/A _1098_/C _1098_/D VGND VGND VPWR VPWR _1102_/Y sky130_fd_sc_hd__o21bai_1
X_1033_ _1834_/Q VGND VGND VPWR VPWR _1421_/B sky130_fd_sc_hd__buf_2
XFILLER_21_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1797_ _1816_/Q _1797_/D VGND VGND VPWR VPWR _1797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1720_ _1760_/Q _1760_/D _1716_/X _1719_/X VGND VGND VPWR VPWR _1840_/D sky130_fd_sc_hd__a31o_1
X_1651_ _1675_/A _1651_/B VGND VGND VPWR VPWR _1652_/A sky130_fd_sc_hd__and2_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1582_ _1817_/Q _1803_/Q VGND VGND VPWR VPWR _1582_/X sky130_fd_sc_hd__and2b_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1016_ _1822_/Q VGND VGND VPWR VPWR _1388_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1849_ _1816_/Q _1849_/D VGND VGND VPWR VPWR _1849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1634_ _1632_/X _1634_/B VGND VGND VPWR VPWR _1635_/A sky130_fd_sc_hd__and2b_1
X_1703_ _1796_/Q _1798_/Q _1703_/C VGND VGND VPWR VPWR _1703_/X sky130_fd_sc_hd__and3_1
XFILLER_39_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1496_ _1493_/X _1494_/X _1500_/A VGND VGND VPWR VPWR _1496_/Y sky130_fd_sc_hd__o21ai_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1565_ _1647_/A input5/X VGND VGND VPWR VPWR _1566_/A sky130_fd_sc_hd__and2_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1350_ _1350_/A _1350_/B _1350_/C VGND VGND VPWR VPWR _1398_/B sky130_fd_sc_hd__and3_1
X_1281_ _1281_/A _1223_/B VGND VGND VPWR VPWR _1283_/A sky130_fd_sc_hd__or2b_1
X_0996_ _0998_/B VGND VGND VPWR VPWR _0996_/Y sky130_fd_sc_hd__inv_2
X_1617_ _1628_/A _1617_/B VGND VGND VPWR VPWR _1617_/Y sky130_fd_sc_hd__nand2_1
XFILLER_54_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1548_ _1548_/A VGND VGND VPWR VPWR _1825_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1479_ _1776_/Q _1780_/Q _1708_/B VGND VGND VPWR VPWR _1498_/B sky130_fd_sc_hd__mux2_1
XFILLER_42_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1402_ _1402_/A _1402_/B _1402_/C VGND VGND VPWR VPWR _1403_/C sky130_fd_sc_hd__nand3_1
XFILLER_5_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput4 rst VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__buf_2
X_1333_ _1318_/B _1319_/A _1320_/B _1320_/A VGND VGND VPWR VPWR _1368_/A sky130_fd_sc_hd__o22a_1
X_1264_ _1246_/X _1318_/A _1264_/C VGND VGND VPWR VPWR _1318_/B sky130_fd_sc_hd__nand3b_1
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1195_ _1195_/A VGND VGND VPWR VPWR _1195_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_24_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0979_ _1282_/B _0979_/B VGND VGND VPWR VPWR _1028_/B sky130_fd_sc_hd__nand2_1
XFILLER_59_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0902_ _1827_/Q _0921_/A _0921_/B _0900_/Y _1155_/A VGND VGND VPWR VPWR _0902_/X
+ sky130_fd_sc_hd__a41o_1
X_1247_ _1823_/Q VGND VGND VPWR VPWR _1347_/A sky130_fd_sc_hd__clkbuf_2
X_1316_ _1315_/A _1295_/A _1315_/C VGND VGND VPWR VPWR _1317_/B sky130_fd_sc_hd__o21a_1
X_1178_ _1178_/A _1277_/C VGND VGND VPWR VPWR _1178_/Y sky130_fd_sc_hd__nand2_1
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1101_ _1101_/A _1101_/B _1101_/C _1101_/D VGND VGND VPWR VPWR _1101_/X sky130_fd_sc_hd__or4_1
X_1032_ _1069_/A VGND VGND VPWR VPWR _1061_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1796_ _1816_/Q _1796_/D VGND VGND VPWR VPWR _1796_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1581_ _1581_/A VGND VGND VPWR VPWR _1765_/D sky130_fd_sc_hd__clkbuf_1
X_1650_ _1778_/Q _1808_/Q _1650_/S VGND VGND VPWR VPWR _1651_/B sky130_fd_sc_hd__mux2_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1015_ _0988_/A _0988_/B _0972_/B VGND VGND VPWR VPWR _1057_/A sky130_fd_sc_hd__o21ai_1
XFILLER_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1848_ _1816_/Q _1848_/D VGND VGND VPWR VPWR _1848_/Q sky130_fd_sc_hd__dfxtp_1
X_1779_ _1816_/Q _1779_/D VGND VGND VPWR VPWR _1779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1633_ _1596_/A _1630_/X _1631_/Y _1773_/Q VGND VGND VPWR VPWR _1634_/B sky130_fd_sc_hd__a31o_1
X_1564_ _1679_/A VGND VGND VPWR VPWR _1647_/A sky130_fd_sc_hd__clkbuf_2
X_1702_ _1800_/Q _1799_/Q _1801_/Q _1802_/Q VGND VGND VPWR VPWR _1703_/C sky130_fd_sc_hd__and4_1
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1495_ _1495_/A _1495_/B VGND VGND VPWR VPWR _1500_/A sky130_fd_sc_hd__or2_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1280_ _1195_/X _1320_/A _1268_/Y _1279_/X _1210_/X VGND VGND VPWR VPWR _1280_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0995_ _0995_/A _0995_/B VGND VGND VPWR VPWR _0998_/B sky130_fd_sc_hd__or2_1
X_1547_ _1547_/A _1549_/B VGND VGND VPWR VPWR _1548_/A sky130_fd_sc_hd__and2_1
X_1616_ _1616_/A _1616_/B VGND VGND VPWR VPWR _1617_/B sky130_fd_sc_hd__xnor2_1
XFILLER_5_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1478_ _1835_/Q VGND VGND VPWR VPWR _1708_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_54_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1401_ _1402_/A _1402_/B _1402_/C VGND VGND VPWR VPWR _1403_/B sky130_fd_sc_hd__a21o_1
XFILLER_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1194_ _1194_/A _1194_/B _1287_/B VGND VGND VPWR VPWR _1194_/X sky130_fd_sc_hd__and3_1
X_1332_ _1447_/A _1332_/B VGND VGND VPWR VPWR _1332_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_36_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1263_ _1263_/A _1263_/B _1263_/C VGND VGND VPWR VPWR _1264_/C sky130_fd_sc_hd__or3_1
Xinput5 select VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__clkbuf_1
XFILLER_51_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0978_ _1348_/C VGND VGND VPWR VPWR _1282_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0901_ _1826_/Q VGND VGND VPWR VPWR _1155_/A sky130_fd_sc_hd__clkinv_2
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1315_ _1315_/A _1426_/C _1315_/C VGND VGND VPWR VPWR _1317_/A sky130_fd_sc_hd__nor3_1
XFILLER_64_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1177_ _1178_/A _1277_/C VGND VGND VPWR VPWR _1208_/B sky130_fd_sc_hd__or2_1
X_1246_ _1246_/A _1246_/B _1263_/B VGND VGND VPWR VPWR _1246_/X sky130_fd_sc_hd__or3_1
XFILLER_24_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1100_ _1100_/A _1101_/D _1100_/C VGND VGND VPWR VPWR _1100_/X sky130_fd_sc_hd__or3_1
X_1031_ _1086_/A _1039_/A _1085_/B _0992_/A _1030_/Y VGND VGND VPWR VPWR _1069_/A
+ sky130_fd_sc_hd__a311oi_4
XFILLER_38_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1795_ _1816_/Q _1795_/D VGND VGND VPWR VPWR _1795_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1229_ _1205_/A _1392_/B _1228_/Y _1257_/A VGND VGND VPWR VPWR _1230_/B sky130_fd_sc_hd__o22a_1
XFILLER_44_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1580_ _1764_/Q _1725_/B VGND VGND VPWR VPWR _1581_/A sky130_fd_sc_hd__and2_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1014_ _1388_/A _1205_/A VGND VGND VPWR VPWR _1060_/A sky130_fd_sc_hd__nand2_1
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1847_ _1816_/Q _1847_/D VGND VGND VPWR VPWR _1847_/Q sky130_fd_sc_hd__dfxtp_1
X_1778_ _1816_/Q _1778_/D VGND VGND VPWR VPWR _1778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1701_ _1816_/Q _1708_/A VGND VGND VPWR VPWR _1816_/D sky130_fd_sc_hd__nor2_1
XFILLER_16_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1632_ _1773_/Q _1609_/C _1630_/X _1631_/Y input4/X VGND VGND VPWR VPWR _1632_/X
+ sky130_fd_sc_hd__a41o_1
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1494_ _1495_/A _1495_/B VGND VGND VPWR VPWR _1494_/X sky130_fd_sc_hd__and2_2
X_1563_ _1693_/A VGND VGND VPWR VPWR _1679_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_58_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0994_ _1393_/B VGND VGND VPWR VPWR _1112_/A sky130_fd_sc_hd__clkbuf_2
X_1546_ _1546_/A VGND VGND VPWR VPWR _1824_/D sky130_fd_sc_hd__clkbuf_1
X_1615_ _1769_/Q _1609_/B _1607_/X VGND VGND VPWR VPWR _1616_/B sky130_fd_sc_hd__a21oi_1
X_1477_ _1793_/Q _0884_/A _1468_/X _1773_/Q VGND VGND VPWR VPWR _1811_/D sky130_fd_sc_hd__a22o_1
XFILLER_5_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1400_ _1400_/A _1400_/B VGND VGND VPWR VPWR _1402_/C sky130_fd_sc_hd__xnor2_1
X_1331_ _1393_/A _1290_/B _1322_/Y VGND VGND VPWR VPWR _1332_/B sky130_fd_sc_hd__a21oi_1
XFILLER_36_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1262_ _1263_/A _1263_/B _1263_/C VGND VGND VPWR VPWR _1318_/A sky130_fd_sc_hd__o21ai_2
X_1193_ _1193_/A VGND VGND VPWR VPWR _1193_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_51_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0977_ _0968_/B _0968_/C _0953_/Y _0954_/Y _0976_/Y VGND VGND VPWR VPWR _0980_/A
+ sky130_fd_sc_hd__o311a_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1529_ _1529_/A VGND VGND VPWR VPWR _1832_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_19_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0900_ _1829_/Q _1828_/Q VGND VGND VPWR VPWR _0900_/Y sky130_fd_sc_hd__nor2_1
XFILLER_33_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1314_ _1314_/A _1314_/B VGND VGND VPWR VPWR _1315_/C sky130_fd_sc_hd__or2_1
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1176_ _1272_/B _1273_/A VGND VGND VPWR VPWR _1277_/C sky130_fd_sc_hd__nand2_1
X_1245_ _1245_/A _1246_/B _1263_/B VGND VGND VPWR VPWR _1268_/A sky130_fd_sc_hd__or3_1
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1030_ _1387_/B _1093_/A VGND VGND VPWR VPWR _1030_/Y sky130_fd_sc_hd__nor2_1
XFILLER_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1794_ _1794_/D _1551_/Y VGND VGND VPWR VPWR _1794_/Q sky130_fd_sc_hd__dlxtn_1
X_1228_ _1228_/A VGND VGND VPWR VPWR _1228_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1159_ _1181_/A VGND VGND VPWR VPWR _1315_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1013_ _1387_/A VGND VGND VPWR VPWR _1205_/A sky130_fd_sc_hd__clkinv_2
XFILLER_34_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1846_ _1816_/Q _1846_/D VGND VGND VPWR VPWR _1846_/Q sky130_fd_sc_hd__dfxtp_1
X_1777_ _1816_/Q _1777_/D VGND VGND VPWR VPWR _1777_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1631_ _1547_/A _1625_/X _1620_/B VGND VGND VPWR VPWR _1631_/Y sky130_fd_sc_hd__o21ai_1
X_1700_ _1853_/Q _1851_/D _1696_/X _1699_/X VGND VGND VPWR VPWR _1803_/D sky130_fd_sc_hd__a31o_1
X_1562_ _1562_/A VGND VGND VPWR VPWR _1757_/D sky130_fd_sc_hd__clkbuf_1
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1493_ _1498_/C VGND VGND VPWR VPWR _1493_/X sky130_fd_sc_hd__buf_2
XFILLER_39_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1829_ _1829_/D _1666_/A VGND VGND VPWR VPWR _1829_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0993_ _1282_/B VGND VGND VPWR VPWR _1393_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_44_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1614_ _1614_/A _1613_/Y VGND VGND VPWR VPWR _1616_/A sky130_fd_sc_hd__or2b_1
X_1545_ _1545_/A _1549_/B VGND VGND VPWR VPWR _1546_/A sky130_fd_sc_hd__and2_1
X_1476_ _1792_/Q _0884_/A _1468_/X _1547_/A VGND VGND VPWR VPWR _1810_/D sky130_fd_sc_hd__a22o_1
XFILLER_54_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1330_ _1330_/A VGND VGND VPWR VPWR _1447_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1261_ _1313_/B _1261_/B VGND VGND VPWR VPWR _1263_/C sky130_fd_sc_hd__and2_1
XFILLER_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1192_ _1192_/A VGND VGND VPWR VPWR _1193_/A sky130_fd_sc_hd__clkbuf_2
X_0976_ _1348_/C VGND VGND VPWR VPWR _0976_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1528_ _1545_/A _1530_/B _1532_/C VGND VGND VPWR VPWR _1529_/A sky130_fd_sc_hd__and3_1
X_1459_ _1786_/Q _1818_/D _1805_/D _1534_/A VGND VGND VPWR VPWR _1812_/D sky130_fd_sc_hd__a22o_1
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1244_ _1244_/A _1244_/B _1287_/B VGND VGND VPWR VPWR _1244_/X sky130_fd_sc_hd__and3_1
X_1313_ _1313_/A _1313_/B _1313_/C VGND VGND VPWR VPWR _1314_/B sky130_fd_sc_hd__and3_1
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR _1839_/CLK sky130_fd_sc_hd__clkbuf_2
X_1175_ _1421_/A _1392_/B VGND VGND VPWR VPWR _1273_/A sky130_fd_sc_hd__nand2_1
X_0959_ _1830_/Q VGND VGND VPWR VPWR _1348_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_32_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1793_ _1793_/D _1551_/Y VGND VGND VPWR VPWR _1793_/Q sky130_fd_sc_hd__dlxtn_1
X_1227_ _1257_/A _1304_/B _1387_/A _1228_/A VGND VGND VPWR VPWR _1257_/B sky130_fd_sc_hd__and4b_1
X_1158_ _1158_/A _1335_/A VGND VGND VPWR VPWR _1181_/A sky130_fd_sc_hd__nand2_1
X_1089_ _1194_/A _1194_/B _0991_/B VGND VGND VPWR VPWR _1089_/X sky130_fd_sc_hd__a21o_1
XFILLER_52_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1012_ _1821_/Q VGND VGND VPWR VPWR _1387_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_34_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1845_ _1816_/Q _1845_/D VGND VGND VPWR VPWR _1845_/Q sky130_fd_sc_hd__dfxtp_1
X_1776_ _1816_/Q _1776_/D VGND VGND VPWR VPWR _1776_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1630_ _1772_/Q _1771_/Q _1625_/X _1624_/B VGND VGND VPWR VPWR _1630_/X sky130_fd_sc_hd__a31o_1
XFILLER_3_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1492_ _1505_/A _1498_/C _1504_/A _1491_/X VGND VGND VPWR VPWR _1492_/X sky130_fd_sc_hd__a31o_1
X_1561_ _1817_/Q _1575_/B VGND VGND VPWR VPWR _1562_/A sky130_fd_sc_hd__and2_1
XFILLER_39_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1828_ _1828_/D _1666_/A VGND VGND VPWR VPWR _1828_/Q sky130_fd_sc_hd__dlxtn_1
X_1759_ _1816_/Q _1759_/D VGND VGND VPWR VPWR _1759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0992_ _0992_/A _0992_/B VGND VGND VPWR VPWR _1086_/A sky130_fd_sc_hd__nor2_2
XFILLER_44_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1544_ _1544_/A VGND VGND VPWR VPWR _1823_/D sky130_fd_sc_hd__clkbuf_1
X_1613_ _1613_/A _1613_/B VGND VGND VPWR VPWR _1613_/Y sky130_fd_sc_hd__nand2_1
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1475_ _1772_/Q VGND VGND VPWR VPWR _1547_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_27_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1260_ _1260_/A _1260_/B VGND VGND VPWR VPWR _1261_/B sky130_fd_sc_hd__nand2_1
X_1191_ _1191_/A VGND VGND VPWR VPWR _1787_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_36_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0975_ _0999_/A _0997_/A _0997_/B _0974_/X VGND VGND VPWR VPWR _0981_/A sky130_fd_sc_hd__a31oi_1
XFILLER_32_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1527_ _1527_/A VGND VGND VPWR VPWR _1831_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1389_ _1388_/A _1826_/Q _1426_/A _1388_/C VGND VGND VPWR VPWR _1389_/X sky130_fd_sc_hd__a22o_1
X_1458_ _1806_/D VGND VGND VPWR VPWR _1534_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1174_ _1197_/A _1198_/B VGND VGND VPWR VPWR _1272_/B sky130_fd_sc_hd__nand2_1
X_1312_ _1313_/A _1313_/B _1313_/C VGND VGND VPWR VPWR _1314_/A sky130_fd_sc_hd__a21oi_1
X_1243_ _1807_/Q _1806_/Q _1223_/Y _1242_/X _1217_/X VGND VGND VPWR VPWR _1789_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0958_ _1830_/Q _0932_/X _0941_/X _0985_/A _0907_/B VGND VGND VPWR VPWR _1244_/A
+ sky130_fd_sc_hd__a311oi_4
X_0889_ _1832_/Q VGND VGND VPWR VPWR _1341_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_20_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1792_ _1792_/D _1551_/Y VGND VGND VPWR VPWR _1792_/Q sky130_fd_sc_hd__dlxtn_1
X_1226_ _1819_/Q _1393_/B _1253_/C VGND VGND VPWR VPWR _1228_/A sky130_fd_sc_hd__a21o_1
X_1157_ _1151_/Y _1155_/Y _1179_/B VGND VGND VPWR VPWR _1157_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_37_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1088_ _1062_/S _1086_/X _1087_/X _1426_/B VGND VGND VPWR VPWR _1142_/A sky130_fd_sc_hd__a211oi_2
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR _1837_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1011_ _1339_/A VGND VGND VPWR VPWR _1388_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_34_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1844_ _1816_/Q _1844_/D VGND VGND VPWR VPWR _1844_/Q sky130_fd_sc_hd__dfxtp_1
X_1775_ _1816_/Q _1775_/D VGND VGND VPWR VPWR _1775_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1209_ _1276_/A _1209_/B VGND VGND VPWR VPWR _1209_/X sky130_fd_sc_hd__xor2_1
XFILLER_25_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1560_ _1690_/A VGND VGND VPWR VPWR _1575_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1491_ _1495_/A VGND VGND VPWR VPWR _1491_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_47_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1827_ _1827_/D _1666_/A VGND VGND VPWR VPWR _1827_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_22_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1689_ _1689_/A VGND VGND VPWR VPWR _1801_/D sky130_fd_sc_hd__clkbuf_1
X_1758_ _1816_/Q _1758_/D VGND VGND VPWR VPWR _1758_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0991_ _1388_/C _0991_/B VGND VGND VPWR VPWR _0992_/B sky130_fd_sc_hd__and2_1
X_1543_ _1613_/A _1549_/B VGND VGND VPWR VPWR _1544_/A sky130_fd_sc_hd__and2_1
X_1474_ _1791_/Q _0884_/A _1468_/X _1545_/A VGND VGND VPWR VPWR _1809_/D sky130_fd_sc_hd__a22o_1
X_1612_ _1770_/Q _1613_/B VGND VGND VPWR VPWR _1614_/A sky130_fd_sc_hd__nor2_1
XFILLER_39_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1190_ _1735_/B _1190_/B _1190_/C VGND VGND VPWR VPWR _1191_/A sky130_fd_sc_hd__and3_1
XFILLER_36_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0974_ _0995_/A _0995_/B _1204_/B VGND VGND VPWR VPWR _0974_/X sky130_fd_sc_hd__o21a_1
XFILLER_32_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1526_ _1613_/A _1530_/B _1532_/C VGND VGND VPWR VPWR _1527_/A sky130_fd_sc_hd__and3_1
X_1457_ _1457_/A VGND VGND VPWR VPWR _1794_/D sky130_fd_sc_hd__clkbuf_1
X_1388_ _1388_/A _1388_/B _1388_/C VGND VGND VPWR VPWR _1388_/X sky130_fd_sc_hd__and3_1
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1311_ _1360_/B _1311_/B VGND VGND VPWR VPWR _1313_/C sky130_fd_sc_hd__nand2_1
XFILLER_64_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1242_ _1008_/S _1287_/B _1241_/X VGND VGND VPWR VPWR _1242_/X sky130_fd_sc_hd__a21o_1
X_1173_ _1192_/A VGND VGND VPWR VPWR _1173_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_2_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0957_ _0961_/B _0961_/C _0968_/B _0968_/C VGND VGND VPWR VPWR _0995_/A sky130_fd_sc_hd__o2bb2a_1
X_0888_ _1554_/A _1556_/A VGND VGND VPWR VPWR _1805_/D sky130_fd_sc_hd__nor2_1
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1509_ _1498_/C _1504_/A _1512_/A VGND VGND VPWR VPWR _1511_/A sky130_fd_sc_hd__mux2_1
XFILLER_55_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1791_ _1791_/D _1551_/Y VGND VGND VPWR VPWR _1791_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1087_ _1061_/A _1061_/B _0991_/B VGND VGND VPWR VPWR _1087_/X sky130_fd_sc_hd__o21a_1
X_1225_ _1225_/A _1225_/B VGND VGND VPWR VPWR _1257_/A sky130_fd_sc_hd__nor2_1
X_1156_ _1806_/Q VGND VGND VPWR VPWR _1179_/B sky130_fd_sc_hd__inv_2
XFILLER_25_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1010_ _1018_/A VGND VGND VPWR VPWR _1339_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1843_ _1816_/Q _1843_/D VGND VGND VPWR VPWR _1843_/Q sky130_fd_sc_hd__dfxtp_1
X_1774_ _1816_/Q _1774_/D VGND VGND VPWR VPWR _1774_/Q sky130_fd_sc_hd__dfxtp_1
X_1208_ _1273_/A _1208_/B VGND VGND VPWR VPWR _1209_/B sky130_fd_sc_hd__nand2_1
XFILLER_27_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1139_ _1121_/X _1126_/X _1138_/X _1110_/X _1249_/B VGND VGND VPWR VPWR _1139_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1490_ _1775_/Q _1779_/Q _1835_/Q VGND VGND VPWR VPWR _1495_/A sky130_fd_sc_hd__mux2_1
XFILLER_54_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1826_ _1826_/D _0880_/X VGND VGND VPWR VPWR _1826_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1688_ _1688_/A _1800_/Q VGND VGND VPWR VPWR _1689_/A sky130_fd_sc_hd__and2_1
X_1757_ _1816_/Q _1757_/D VGND VGND VPWR VPWR _1757_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0990_ _1388_/C _0991_/B VGND VGND VPWR VPWR _0992_/A sky130_fd_sc_hd__nor2_2
X_1611_ _1541_/A _1609_/X _1610_/X VGND VGND VPWR VPWR _1769_/D sky130_fd_sc_hd__o21ba_1
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1542_ _1542_/A VGND VGND VPWR VPWR _1822_/D sky130_fd_sc_hd__clkbuf_1
X_1473_ _1771_/Q VGND VGND VPWR VPWR _1545_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_39_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1809_ _1809_/D _1667_/B VGND VGND VPWR VPWR _1809_/Q sky130_fd_sc_hd__dlxtn_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0973_ _1020_/A _1004_/A _1004_/B _1007_/A VGND VGND VPWR VPWR _0997_/B sky130_fd_sc_hd__a31o_1
X_1387_ _1387_/A _1387_/B VGND VGND VPWR VPWR _1391_/A sky130_fd_sc_hd__nand2_1
X_1525_ _1525_/A VGND VGND VPWR VPWR _1830_/D sky130_fd_sc_hd__clkbuf_1
X_1456_ _1456_/A _1456_/B _1456_/C VGND VGND VPWR VPWR _1457_/A sky130_fd_sc_hd__and3_1
XFILLER_35_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1310_ _1310_/A _1310_/B VGND VGND VPWR VPWR _1311_/B sky130_fd_sc_hd__or2_1
X_1241_ _1195_/A _1238_/X _1240_/Y _1210_/A _1173_/X VGND VGND VPWR VPWR _1241_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1172_ _1807_/Q _1806_/Q VGND VGND VPWR VPWR _1192_/A sky130_fd_sc_hd__nor2_1
XFILLER_2_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0956_ _0956_/A VGND VGND VPWR VPWR _1204_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_32_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_0887_ _0887_/A VGND VGND VPWR VPWR _0887_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1439_ _1407_/A _1437_/Y _1438_/X VGND VGND VPWR VPWR _1442_/A sky130_fd_sc_hd__a21o_1
X_1508_ _1493_/X _1494_/X _1503_/X _1505_/A _1507_/Y VGND VGND VPWR VPWR _1508_/Y
+ sky130_fd_sc_hd__o221ai_4
XFILLER_62_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1790_ _1790_/D _1551_/Y VGND VGND VPWR VPWR _1790_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_14_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1224_ _1341_/C _1393_/B VGND VGND VPWR VPWR _1225_/B sky130_fd_sc_hd__nand2_1
XFILLER_37_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1086_ _1086_/A _1086_/B VGND VGND VPWR VPWR _1086_/X sky130_fd_sc_hd__xor2_2
XFILLER_52_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1155_ _1155_/A _1155_/B VGND VGND VPWR VPWR _1155_/Y sky130_fd_sc_hd__nand2_1
XFILLER_16_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0939_ _0966_/A _1823_/Q VGND VGND VPWR VPWR _0968_/A sky130_fd_sc_hd__nor2_1
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1773_ _1816_/Q _1773_/D VGND VGND VPWR VPWR _1773_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_8_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1842_ _1816_/Q _1842_/D VGND VGND VPWR VPWR _1842_/Q sky130_fd_sc_hd__dfxtp_1
X_1207_ _1207_/A VGND VGND VPWR VPWR _1276_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1069_ _1069_/A _1069_/B _1069_/C _1201_/A VGND VGND VPWR VPWR _1070_/B sky130_fd_sc_hd__or4b_1
X_1138_ _1420_/B _1126_/B _1126_/C _1136_/X _1137_/X VGND VGND VPWR VPWR _1138_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_43_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1825_ _1825_/D _0880_/X VGND VGND VPWR VPWR _1825_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_30_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1756_ _1756_/A VGND VGND VPWR VPWR _1857_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1687_ _1687_/A VGND VGND VPWR VPWR _1800_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1610_ _1541_/A _1609_/X _1711_/S VGND VGND VPWR VPWR _1610_/X sky130_fd_sc_hd__a21o_1
XFILLER_8_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1541_ _1541_/A _1549_/B VGND VGND VPWR VPWR _1542_/A sky130_fd_sc_hd__and2_1
X_1472_ _1790_/Q _0884_/A _1468_/X _1613_/A VGND VGND VPWR VPWR _1808_/D sky130_fd_sc_hd__a22o_1
XFILLER_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1739_ _1845_/Q _1848_/Q _1847_/Q VGND VGND VPWR VPWR _1739_/X sky130_fd_sc_hd__and3_1
X_1808_ _1808_/D _1667_/B VGND VGND VPWR VPWR _1808_/Q sky130_fd_sc_hd__dlxtn_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0972_ _1018_/A _0972_/B VGND VGND VPWR VPWR _1007_/A sky130_fd_sc_hd__nand2_1
XFILLER_32_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1524_ _1541_/A _1530_/B _1532_/C VGND VGND VPWR VPWR _1525_/A sky130_fd_sc_hd__and3_1
X_1386_ _1386_/A _1386_/B VGND VGND VPWR VPWR _1403_/A sky130_fd_sc_hd__xor2_1
X_1455_ _1376_/A _1155_/B _1454_/X _1806_/Q _1807_/Q VGND VGND VPWR VPWR _1456_/C
+ sky130_fd_sc_hd__a2111o_1
XFILLER_42_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1171_ _1171_/A VGND VGND VPWR VPWR _1287_/B sky130_fd_sc_hd__clkbuf_2
X_1240_ _1281_/A _1240_/B VGND VGND VPWR VPWR _1240_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0955_ _0968_/B _0968_/C _0953_/Y _0954_/Y VGND VGND VPWR VPWR _0979_/B sky130_fd_sc_hd__o31ai_2
X_0886_ _1838_/Q _1665_/A _1837_/Q VGND VGND VPWR VPWR _0887_/A sky130_fd_sc_hd__and3b_1
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1507_ _1507_/A VGND VGND VPWR VPWR _1507_/Y sky130_fd_sc_hd__inv_2
XFILLER_55_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1438_ _1438_/A _1438_/B VGND VGND VPWR VPWR _1438_/X sky130_fd_sc_hd__and2_1
X_1369_ _1368_/A _1368_/B _1195_/A VGND VGND VPWR VPWR _1369_/X sky130_fd_sc_hd__a21bo_1
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1154_ _1111_/X _1139_/X _1151_/Y _1153_/X VGND VGND VPWR VPWR _1154_/X sky130_fd_sc_hd__a211o_1
X_1223_ _1281_/A _1223_/B VGND VGND VPWR VPWR _1223_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1085_ _1085_/A _1085_/B VGND VGND VPWR VPWR _1086_/B sky130_fd_sc_hd__nand2_1
XFILLER_37_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0938_ _0961_/B _0961_/C _1350_/B VGND VGND VPWR VPWR _0962_/B sky130_fd_sc_hd__a21o_1
XFILLER_57_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1772_ _1816_/Q _1772_/D VGND VGND VPWR VPWR _1772_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1841_ _1816_/Q _1841_/D VGND VGND VPWR VPWR _1841_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1137_ _1137_/A _1178_/A VGND VGND VPWR VPWR _1137_/X sky130_fd_sc_hd__and2_1
X_1206_ _1206_/A _1206_/B VGND VGND VPWR VPWR _1207_/A sky130_fd_sc_hd__nor2_1
XFILLER_25_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1068_ _1158_/A _1422_/A VGND VGND VPWR VPWR _1201_/A sky130_fd_sc_hd__nand2_1
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1824_ _1824_/D _0880_/X VGND VGND VPWR VPWR _1824_/Q sky130_fd_sc_hd__dlxtn_1
X_1755_ _1755_/A _1856_/Q VGND VGND VPWR VPWR _1756_/A sky130_fd_sc_hd__and2_1
X_1686_ _1688_/A _1799_/Q VGND VGND VPWR VPWR _1687_/A sky130_fd_sc_hd__and2_1
XFILLER_57_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1540_ _1540_/A VGND VGND VPWR VPWR _1549_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1471_ _1770_/Q VGND VGND VPWR VPWR _1613_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1807_ _1807_/D _0887_/X VGND VGND VPWR VPWR _1807_/Q sky130_fd_sc_hd__dlxtp_1
XFILLER_49_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1669_ _1665_/X _1666_/Y _1667_/Y _1668_/X _1783_/Q VGND VGND VPWR VPWR _1783_/D
+ sky130_fd_sc_hd__a32o_1
X_1738_ _1842_/Q _1841_/Q _1844_/Q _1843_/Q VGND VGND VPWR VPWR _1738_/X sky130_fd_sc_hd__or4_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0971_ _1822_/Q VGND VGND VPWR VPWR _0972_/B sky130_fd_sc_hd__inv_2
XFILLER_32_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1523_ _1523_/A VGND VGND VPWR VPWR _1532_/C sky130_fd_sc_hd__clkbuf_1
X_1454_ _1376_/A _1155_/B _1379_/B VGND VGND VPWR VPWR _1454_/X sky130_fd_sc_hd__o21a_1
XFILLER_55_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1385_ _1385_/A _1384_/X VGND VGND VPWR VPWR _1386_/B sky130_fd_sc_hd__or2b_1
XFILLER_27_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1170_ _1183_/A _1179_/B VGND VGND VPWR VPWR _1171_/A sky130_fd_sc_hd__nor2_1
XFILLER_37_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0954_ _0968_/B _0968_/C _0951_/B VGND VGND VPWR VPWR _0954_/Y sky130_fd_sc_hd__o21ai_1
X_0885_ _1836_/Q VGND VGND VPWR VPWR _1665_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1437_ _1437_/A VGND VGND VPWR VPWR _1437_/Y sky130_fd_sc_hd__inv_2
X_1506_ _1485_/A _1493_/X _1503_/X _1505_/X VGND VGND VPWR VPWR _1506_/X sky130_fd_sc_hd__o31a_2
XFILLER_55_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1299_ _1334_/A _1341_/B _1299_/C _1300_/A VGND VGND VPWR VPWR _1334_/B sky130_fd_sc_hd__and4b_1
X_1368_ _1368_/A _1368_/B VGND VGND VPWR VPWR _1409_/B sky130_fd_sc_hd__nor2_1
XFILLER_11_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1084_ _1084_/A _1084_/B VGND VGND VPWR VPWR _1084_/Y sky130_fd_sc_hd__xnor2_1
X_1153_ _1290_/B _1106_/X _1145_/X _1422_/B _1152_/X VGND VGND VPWR VPWR _1153_/X
+ sky130_fd_sc_hd__a221o_1
X_1222_ _1222_/A _1345_/A VGND VGND VPWR VPWR _1223_/B sky130_fd_sc_hd__or2b_1
XFILLER_60_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0937_ _0937_/A VGND VGND VPWR VPWR _1350_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_9_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1840_ _1816_/Q _1840_/D VGND VGND VPWR VPWR _1840_/Q sky130_fd_sc_hd__dfxtp_1
X_1771_ _1816_/Q _1771_/D VGND VGND VPWR VPWR _1771_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1205_ _1205_/A _1205_/B VGND VGND VPWR VPWR _1206_/B sky130_fd_sc_hd__nor2_1
X_1067_ _1158_/A _1422_/A VGND VGND VPWR VPWR _1069_/B sky130_fd_sc_hd__nor2_1
X_1136_ _1197_/A _1124_/S _1178_/A _1137_/A _1135_/X VGND VGND VPWR VPWR _1136_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_40_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1823_ _1823_/D _0880_/X VGND VGND VPWR VPWR _1823_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_15_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1754_ _1754_/A VGND VGND VPWR VPWR _1856_/D sky130_fd_sc_hd__clkbuf_1
X_1685_ _1685_/A VGND VGND VPWR VPWR _1799_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_57_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1119_ _1100_/X _1103_/X _1116_/X _1117_/Y _1376_/B VGND VGND VPWR VPWR _1119_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1470_ _1789_/Q _1818_/D _1468_/X _1541_/A VGND VGND VPWR VPWR _1815_/D sky130_fd_sc_hd__a22o_1
XFILLER_8_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1806_ _1806_/D _0887_/X VGND VGND VPWR VPWR _1806_/Q sky130_fd_sc_hd__dlxtp_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1668_ _1679_/A _1668_/B _1668_/C VGND VGND VPWR VPWR _1668_/X sky130_fd_sc_hd__and3_1
X_1599_ _1755_/A VGND VGND VPWR VPWR _1599_/X sky130_fd_sc_hd__clkbuf_2
X_1737_ _1846_/Q _1845_/Q _1848_/Q _1847_/Q VGND VGND VPWR VPWR _1737_/X sky130_fd_sc_hd__or4_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0970_ _1004_/A _1004_/B _1020_/A VGND VGND VPWR VPWR _0997_/A sky130_fd_sc_hd__a21o_1
XFILLER_32_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1522_ _1522_/A VGND VGND VPWR VPWR _1829_/D sky130_fd_sc_hd__clkbuf_1
X_1453_ _1195_/X _1445_/Y _1452_/X _1173_/X VGND VGND VPWR VPWR _1456_/B sky130_fd_sc_hd__a211o_1
X_1384_ _1180_/A _1833_/Q _1339_/X _1344_/A VGND VGND VPWR VPWR _1384_/X sky130_fd_sc_hd__a211o_1
XFILLER_50_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_0953_ _0953_/A _0953_/B VGND VGND VPWR VPWR _0953_/Y sky130_fd_sc_hd__xnor2_1
X_0884_ _0884_/A VGND VGND VPWR VPWR _1818_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1436_ _1436_/A _1436_/B VGND VGND VPWR VPWR _1443_/A sky130_fd_sc_hd__xnor2_1
X_1367_ _1409_/A _1367_/B VGND VGND VPWR VPWR _1368_/B sky130_fd_sc_hd__or2_1
X_1505_ _1505_/A _1505_/B _1512_/C VGND VGND VPWR VPWR _1505_/X sky130_fd_sc_hd__or3_1
XFILLER_63_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1298_ _1339_/A _1393_/A _1341_/C _1339_/D VGND VGND VPWR VPWR _1300_/A sky130_fd_sc_hd__a22o_1
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1221_ _1821_/Q _1221_/B VGND VGND VPWR VPWR _1345_/A sky130_fd_sc_hd__nand2_2
X_1083_ _1101_/A _1109_/A VGND VGND VPWR VPWR _1084_/B sky130_fd_sc_hd__or2b_1
X_1152_ _1155_/A _1155_/B VGND VGND VPWR VPWR _1152_/X sky130_fd_sc_hd__and2_1
XFILLER_37_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0936_ _0945_/A _0945_/B _0935_/C _1290_/A VGND VGND VPWR VPWR _0961_/C sky130_fd_sc_hd__a31o_1
XFILLER_45_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1419_ _1422_/A _1426_/B _1389_/X _1388_/X _1826_/Q VGND VGND VPWR VPWR _1425_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_28_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1770_ _1816_/Q _1770_/D VGND VGND VPWR VPWR _1770_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1204_ _1422_/A _1204_/B VGND VGND VPWR VPWR _1206_/A sky130_fd_sc_hd__nor2_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1135_ _1100_/X _1103_/X _1134_/Y _1376_/B VGND VGND VPWR VPWR _1135_/X sky130_fd_sc_hd__a211o_1
X_1066_ _1387_/A VGND VGND VPWR VPWR _1422_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_33_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0919_ _0919_/A _0946_/B _0934_/A VGND VGND VPWR VPWR _0920_/B sky130_fd_sc_hd__and3_1
XFILLER_0_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1822_ _1822_/D _0880_/X VGND VGND VPWR VPWR _1822_/Q sky130_fd_sc_hd__dlxtn_1
X_1753_ _1755_/A _1855_/Q VGND VGND VPWR VPWR _1754_/A sky130_fd_sc_hd__and2_1
X_1684_ _1688_/A _1798_/Q VGND VGND VPWR VPWR _1685_/A sky130_fd_sc_hd__and2_1
X_1049_ _1101_/C _1101_/D VGND VGND VPWR VPWR _1084_/A sky130_fd_sc_hd__nor2_1
XFILLER_53_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1118_ _1421_/B VGND VGND VPWR VPWR _1376_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1805_ _1805_/D _1555_/X VGND VGND VPWR VPWR _1805_/Q sky130_fd_sc_hd__dlxtn_1
X_1736_ _1736_/A VGND VGND VPWR VPWR _1848_/D sky130_fd_sc_hd__clkbuf_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1667_ _1849_/Q _1667_/B VGND VGND VPWR VPWR _1667_/Y sky130_fd_sc_hd__nor2_1
X_1598_ _1690_/A VGND VGND VPWR VPWR _1755_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1383_ _1339_/X _1344_/A _1180_/A _1335_/B VGND VGND VPWR VPWR _1385_/A sky130_fd_sc_hd__o211a_1
X_1452_ _1278_/B _1446_/Y _1447_/Y _1451_/X _1210_/A VGND VGND VPWR VPWR _1452_/X
+ sky130_fd_sc_hd__o311a_1
X_1521_ _1603_/A _1532_/B _1523_/A VGND VGND VPWR VPWR _1522_/A sky130_fd_sc_hd__and3_1
XFILLER_35_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1719_ _1717_/X _1718_/X _1840_/Q _1679_/A VGND VGND VPWR VPWR _1719_/X sky130_fd_sc_hd__o211a_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0952_ _0952_/A _0983_/B VGND VGND VPWR VPWR _0953_/B sky130_fd_sc_hd__nor2_1
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0883_ _0883_/A VGND VGND VPWR VPWR _0884_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1504_ _1504_/A _1495_/A VGND VGND VPWR VPWR _1512_/C sky130_fd_sc_hd__or2b_1
XFILLER_55_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1435_ _1400_/A _1400_/B _1399_/A VGND VGND VPWR VPWR _1436_/B sky130_fd_sc_hd__a21oi_1
X_1366_ _1408_/A _1365_/D _1318_/A _1319_/A VGND VGND VPWR VPWR _1367_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1297_ _1339_/A _1393_/A _1341_/C _1339_/D VGND VGND VPWR VPWR _1334_/A sky130_fd_sc_hd__and4_1
XFILLER_11_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1151_ _1422_/B _1145_/X _1149_/X _1155_/B VGND VGND VPWR VPWR _1151_/Y sky130_fd_sc_hd__o22ai_2
X_1220_ _1426_/A _1220_/B VGND VGND VPWR VPWR _1281_/A sky130_fd_sc_hd__xnor2_4
X_1082_ _1116_/A _1082_/B _1082_/C VGND VGND VPWR VPWR _1109_/A sky130_fd_sc_hd__or3_1
XFILLER_52_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0935_ _0945_/A _0945_/B _0935_/C _0935_/D VGND VGND VPWR VPWR _0961_/B sky130_fd_sc_hd__nand4_2
X_1349_ _1345_/B _1347_/Y _1398_/A VGND VGND VPWR VPWR _1350_/C sky130_fd_sc_hd__a21oi_1
X_1418_ _1382_/A _1376_/B _1384_/X _1385_/A VGND VGND VPWR VPWR _1432_/A sky130_fd_sc_hd__a31o_1
XFILLER_51_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1134_ _1158_/A _1421_/A VGND VGND VPWR VPWR _1134_/Y sky130_fd_sc_hd__xnor2_1
X_1203_ _1246_/A _1202_/C _1202_/A VGND VGND VPWR VPWR _1203_/X sky130_fd_sc_hd__a21o_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1065_ _1388_/A VGND VGND VPWR VPWR _1158_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_33_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0918_ _0919_/A _0946_/B _0934_/A VGND VGND VPWR VPWR _0920_/A sky130_fd_sc_hd__a21oi_1
XFILLER_56_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1821_ _1821_/D _0880_/X VGND VGND VPWR VPWR _1821_/Q sky130_fd_sc_hd__dlxtn_2
X_1752_ _1752_/A VGND VGND VPWR VPWR _1855_/D sky130_fd_sc_hd__clkbuf_1
X_1683_ _1683_/A VGND VGND VPWR VPWR _1798_/D sky130_fd_sc_hd__clkbuf_1
X_1117_ _1116_/A _1116_/B _1116_/C VGND VGND VPWR VPWR _1117_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1048_ _1047_/B _1047_/C _1270_/B VGND VGND VPWR VPWR _1101_/D sky130_fd_sc_hd__a21oi_2
XFILLER_53_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1666_ _1666_/A _1672_/S VGND VGND VPWR VPWR _1666_/Y sky130_fd_sc_hd__nand2_1
X_1804_ _1804_/D _1668_/C VGND VGND VPWR VPWR _1804_/Q sky130_fd_sc_hd__dlxtn_1
X_1735_ _1847_/Q _1735_/B VGND VGND VPWR VPWR _1736_/A sky130_fd_sc_hd__and2_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1597_ _1594_/Y _1595_/X _1628_/A VGND VGND VPWR VPWR _1597_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_53_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1520_ _1520_/A VGND VGND VPWR VPWR _1828_/D sky130_fd_sc_hd__clkbuf_1
X_1382_ _1382_/A _1421_/B VGND VGND VPWR VPWR _1386_/A sky130_fd_sc_hd__nand2_1
X_1451_ _1329_/B _1447_/B _1450_/Y _1152_/X VGND VGND VPWR VPWR _1451_/X sky130_fd_sc_hd__a31o_1
XFILLER_23_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1718_ _1758_/Q _1759_/Q _1760_/Q _1761_/Q VGND VGND VPWR VPWR _1718_/X sky130_fd_sc_hd__or4_1
X_1649_ _1679_/A VGND VGND VPWR VPWR _1675_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_58_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0951_ _1348_/D _0951_/B VGND VGND VPWR VPWR _0952_/A sky130_fd_sc_hd__nor2_1
XFILLER_40_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0882_ _1668_/B _1556_/A VGND VGND VPWR VPWR _0883_/A sky130_fd_sc_hd__and2_1
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1503_ _1495_/A _1504_/A VGND VGND VPWR VPWR _1503_/X sky130_fd_sc_hd__and2b_1
X_1434_ _1403_/A _1403_/C _1403_/B VGND VGND VPWR VPWR _1436_/A sky130_fd_sc_hd__a21bo_1
X_1296_ _1350_/A VGND VGND VPWR VPWR _1393_/A sky130_fd_sc_hd__clkbuf_2
X_1365_ _1318_/A _1319_/A _1408_/A _1365_/D VGND VGND VPWR VPWR _1409_/A sky130_fd_sc_hd__and4bb_1
XFILLER_51_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1150_ _1376_/B VGND VGND VPWR VPWR _1155_/B sky130_fd_sc_hd__clkbuf_2
X_1081_ _1101_/A _1101_/B VGND VGND VPWR VPWR _1082_/C sky130_fd_sc_hd__or2_1
XFILLER_60_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0934_ _0934_/A _0934_/B VGND VGND VPWR VPWR _0935_/D sky130_fd_sc_hd__nand2_1
XFILLER_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1417_ _1379_/X _1380_/Y _1217_/X _1416_/X VGND VGND VPWR VPWR _1793_/D sky130_fd_sc_hd__o211a_1
X_1348_ _1823_/Q _1822_/Q _1348_/C _1348_/D VGND VGND VPWR VPWR _1398_/A sky130_fd_sc_hd__and4_1
XFILLER_36_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1279_ _1446_/A _1279_/B VGND VGND VPWR VPWR _1279_/X sky130_fd_sc_hd__xor2_1
XFILLER_51_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1064_ _1194_/A _1194_/B _1205_/A VGND VGND VPWR VPWR _1070_/A sky130_fd_sc_hd__a21o_1
X_1133_ _1133_/A VGND VGND VPWR VPWR _1137_/A sky130_fd_sc_hd__clkbuf_2
X_1202_ _1202_/A _1246_/A _1202_/C VGND VGND VPWR VPWR _1245_/A sky130_fd_sc_hd__nand3_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0917_ _1018_/A _1290_/A VGND VGND VPWR VPWR _0934_/A sky130_fd_sc_hd__nand2_1
XFILLER_56_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1820_ _1820_/D _0880_/X VGND VGND VPWR VPWR _1820_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_30_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1751_ _1755_/A _1854_/Q VGND VGND VPWR VPWR _1752_/A sky130_fd_sc_hd__and2_1
X_1682_ _1688_/A _1797_/Q VGND VGND VPWR VPWR _1683_/A sky130_fd_sc_hd__and2_1
X_1047_ _1270_/B _1047_/B _1047_/C VGND VGND VPWR VPWR _1101_/C sky130_fd_sc_hd__and3_1
X_1116_ _1116_/A _1116_/B _1116_/C VGND VGND VPWR VPWR _1116_/X sky130_fd_sc_hd__or3_1
XFILLER_38_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1803_ _1816_/Q _1803_/D VGND VGND VPWR VPWR _1803_/Q sky130_fd_sc_hd__dfxtp_1
X_1596_ _1596_/A VGND VGND VPWR VPWR _1628_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1665_ _1665_/A _1672_/S VGND VGND VPWR VPWR _1665_/X sky130_fd_sc_hd__or2_1
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1734_ _1734_/A VGND VGND VPWR VPWR _1847_/D sky130_fd_sc_hd__clkbuf_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1450_ _1448_/Y _1446_/Y _1449_/X VGND VGND VPWR VPWR _1450_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1381_ _1381_/A _1361_/X VGND VGND VPWR VPWR _1438_/A sky130_fd_sc_hd__or2b_1
XFILLER_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1579_ _1579_/A VGND VGND VPWR VPWR _1764_/D sky130_fd_sc_hd__clkbuf_1
X_1717_ _1762_/Q _1763_/Q _1764_/Q _1765_/Q VGND VGND VPWR VPWR _1717_/X sky130_fd_sc_hd__or4_1
X_1648_ _1648_/A VGND VGND VPWR VPWR _1777_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0950_ _0950_/A VGND VGND VPWR VPWR _1348_/D sky130_fd_sc_hd__clkbuf_2
X_0881_ _1836_/Q _1837_/Q VGND VGND VPWR VPWR _1556_/A sky130_fd_sc_hd__nor2_1
XFILLER_13_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1433_ _1408_/A _1408_/B _1410_/Y VGND VGND VPWR VPWR _1444_/A sky130_fd_sc_hd__o21ai_1
X_1502_ _1507_/A _1502_/B VGND VGND VPWR VPWR _1502_/Y sky130_fd_sc_hd__nor2_2
XFILLER_55_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1295_ _1295_/A VGND VGND VPWR VPWR _1426_/C sky130_fd_sc_hd__clkbuf_2
X_1364_ _1361_/X _1362_/Y _1314_/A _1317_/A VGND VGND VPWR VPWR _1365_/D sky130_fd_sc_hd__a211o_1
XFILLER_23_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1080_ _1112_/A _1107_/A _1107_/B VGND VGND VPWR VPWR _1101_/B sky130_fd_sc_hd__and3_1
XFILLER_60_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_0933_ _0966_/A _1350_/A VGND VGND VPWR VPWR _0934_/B sky130_fd_sc_hd__nand2_1
X_1347_ _1347_/A _1348_/D VGND VGND VPWR VPWR _1347_/Y sky130_fd_sc_hd__nand2_1
X_1416_ _1195_/X _1409_/X _1410_/Y _1415_/X VGND VGND VPWR VPWR _1416_/X sky130_fd_sc_hd__a31o_1
XFILLER_3_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1278_ _1448_/A _1278_/B VGND VGND VPWR VPWR _1279_/B sky130_fd_sc_hd__nand2_1
XFILLER_24_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1201_ _1201_/A _1201_/B VGND VGND VPWR VPWR _1202_/C sky130_fd_sc_hd__nand2_1
X_1063_ _1205_/B _1114_/B VGND VGND VPWR VPWR _1116_/A sky130_fd_sc_hd__and2_1
X_1132_ _1277_/A VGND VGND VPWR VPWR _1178_/A sky130_fd_sc_hd__clkbuf_2
X_0916_ _1824_/Q VGND VGND VPWR VPWR _1290_/A sky130_fd_sc_hd__inv_2
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1750_ _1750_/A VGND VGND VPWR VPWR _1854_/D sky130_fd_sc_hd__clkbuf_1
X_1681_ _1681_/A VGND VGND VPWR VPWR _1797_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_38_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1115_ _1133_/A _1122_/B _1078_/X VGND VGND VPWR VPWR _1116_/C sky130_fd_sc_hd__o21ai_1
XFILLER_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1046_ _1249_/B VGND VGND VPWR VPWR _1270_/B sky130_fd_sc_hd__clkinv_2
XFILLER_21_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1733_ _1846_/Q _1735_/B VGND VGND VPWR VPWR _1734_/A sky130_fd_sc_hd__and2_1
X_1802_ _1816_/Q _1802_/D VGND VGND VPWR VPWR _1802_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1595_ _1806_/D _1595_/B VGND VGND VPWR VPWR _1595_/X sky130_fd_sc_hd__and2_1
XFILLER_7_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1664_ _1839_/Q _1840_/Q VGND VGND VPWR VPWR _1672_/S sky130_fd_sc_hd__and2b_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1029_ _0985_/B _1008_/S _1028_/X VGND VGND VPWR VPWR _1093_/A sky130_fd_sc_hd__o21ba_1
XFILLER_53_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1380_ _1447_/B _1379_/B _1193_/A VGND VGND VPWR VPWR _1380_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_35_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1716_ _1758_/Q _1761_/Q _1716_/C VGND VGND VPWR VPWR _1716_/X sky130_fd_sc_hd__and3_1
XFILLER_58_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1578_ _1763_/Q _1725_/B VGND VGND VPWR VPWR _1579_/A sky130_fd_sc_hd__and2_1
X_1647_ _1647_/A _1647_/B VGND VGND VPWR VPWR _1648_/A sky130_fd_sc_hd__and2_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0880_ _0880_/A VGND VGND VPWR VPWR _0880_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_13_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1432_ _1432_/A _1432_/B VGND VGND VPWR VPWR _1445_/A sky130_fd_sc_hd__xnor2_2
X_1363_ _1314_/A _1317_/A _1361_/X _1362_/Y VGND VGND VPWR VPWR _1408_/A sky130_fd_sc_hd__o211ai_2
X_1501_ _1491_/X _1505_/A _1500_/Y _1494_/X _1505_/B VGND VGND VPWR VPWR _1502_/B
+ sky130_fd_sc_hd__o221a_1
X_1294_ _1446_/B _1294_/B VGND VGND VPWR VPWR _1294_/X sky130_fd_sc_hd__or2_1
XFILLER_31_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0932_ _0950_/A _0951_/B VGND VGND VPWR VPWR _0932_/X sky130_fd_sc_hd__or2_1
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1346_ _1346_/A _1346_/B VGND VGND VPWR VPWR _1354_/B sky130_fd_sc_hd__nor2_1
X_1415_ _1210_/X _1413_/X _1414_/X _1173_/X VGND VGND VPWR VPWR _1415_/X sky130_fd_sc_hd__a211o_1
XFILLER_28_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1277_ _1277_/A _1277_/B _1277_/C _1277_/D VGND VGND VPWR VPWR _1278_/B sky130_fd_sc_hd__or4_1
XFILLER_36_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1200_ _1201_/A _1201_/B VGND VGND VPWR VPWR _1246_/A sky130_fd_sc_hd__or2_1
X_1062_ _1058_/Y _1060_/Y _1062_/S VGND VGND VPWR VPWR _1114_/B sky130_fd_sc_hd__mux2_2
X_1131_ _1162_/A _1382_/A VGND VGND VPWR VPWR _1277_/A sky130_fd_sc_hd__nor2_1
XFILLER_33_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0915_ _1827_/Q VGND VGND VPWR VPWR _1018_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_33_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1329_ _1329_/A _1329_/B VGND VGND VPWR VPWR _1330_/A sky130_fd_sc_hd__and2_1
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1680_ _1688_/A _1796_/Q VGND VGND VPWR VPWR _1681_/A sky130_fd_sc_hd__and2_1
X_1114_ _1420_/B _1114_/B VGND VGND VPWR VPWR _1116_/B sky130_fd_sc_hd__nor2_1
XFILLER_38_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1045_ _1388_/C VGND VGND VPWR VPWR _1249_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_53_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1732_ _1732_/A VGND VGND VPWR VPWR _1846_/D sky130_fd_sc_hd__clkbuf_1
X_1801_ _1816_/Q _1801_/D VGND VGND VPWR VPWR _1801_/Q sky130_fd_sc_hd__dfxtp_1
X_1663_ _1663_/A VGND VGND VPWR VPWR _1782_/D sky130_fd_sc_hd__clkbuf_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1594_ _1806_/D _1595_/B VGND VGND VPWR VPWR _1594_/Y sky130_fd_sc_hd__nor2_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1028_ _1028_/A _1028_/B _1028_/C VGND VGND VPWR VPWR _1028_/X sky130_fd_sc_hd__and3_1
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1715_ _1762_/Q _1763_/Q _1764_/Q _1765_/Q VGND VGND VPWR VPWR _1716_/C sky130_fd_sc_hd__and4_1
X_1646_ _1777_/Q _1815_/Q _1650_/S VGND VGND VPWR VPWR _1647_/B sky130_fd_sc_hd__mux2_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1577_ _1690_/A VGND VGND VPWR VPWR _1725_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_41_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1500_ _1500_/A VGND VGND VPWR VPWR _1500_/Y sky130_fd_sc_hd__inv_2
X_1431_ _1431_/A _1431_/B VGND VGND VPWR VPWR _1432_/B sky130_fd_sc_hd__xnor2_1
X_1362_ _1381_/A _1361_/C _1361_/A VGND VGND VPWR VPWR _1362_/Y sky130_fd_sc_hd__o21ai_1
X_1293_ _1446_/B _1294_/B VGND VGND VPWR VPWR _1293_/Y sky130_fd_sc_hd__nand2_1
XFILLER_48_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1629_ _1547_/A _1628_/A _1628_/Y _1599_/X VGND VGND VPWR VPWR _1772_/D sky130_fd_sc_hd__o211a_1
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0931_ _0931_/A VGND VGND VPWR VPWR _0951_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_13_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1345_ _1345_/A _1345_/B VGND VGND VPWR VPWR _1354_/A sky130_fd_sc_hd__nor2_1
X_1414_ _1162_/A _1376_/A _0945_/A _0900_/Y _1171_/A VGND VGND VPWR VPWR _1414_/X
+ sky130_fd_sc_hd__o2111a_1
X_1276_ _1276_/A _1281_/A VGND VGND VPWR VPWR _1277_/D sky130_fd_sc_hd__nand2_1
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1130_ _1335_/A VGND VGND VPWR VPWR _1382_/A sky130_fd_sc_hd__clkbuf_2
X_1061_ _1061_/A _1061_/B VGND VGND VPWR VPWR _1062_/S sky130_fd_sc_hd__nor2_1
XFILLER_33_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0914_ _1327_/A _0910_/B _1020_/A VGND VGND VPWR VPWR _0946_/B sky130_fd_sc_hd__a21o_1
X_1328_ _1420_/A _1411_/B VGND VGND VPWR VPWR _1329_/B sky130_fd_sc_hd__nand2_1
X_1259_ _1260_/A _1260_/B VGND VGND VPWR VPWR _1313_/B sky130_fd_sc_hd__or2_1
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1044_ _1047_/B _1047_/C VGND VGND VPWR VPWR _1044_/Y sky130_fd_sc_hd__nand2_1
X_1113_ _1205_/B VGND VGND VPWR VPWR _1420_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1800_ _1816_/Q _1800_/D VGND VGND VPWR VPWR _1800_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1731_ _1845_/Q _1735_/B VGND VGND VPWR VPWR _1732_/A sky130_fd_sc_hd__and2_1
X_1662_ _1803_/Q _1725_/B VGND VGND VPWR VPWR _1663_/A sky130_fd_sc_hd__and2_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1593_ _1807_/D _1624_/B VGND VGND VPWR VPWR _1595_/B sky130_fd_sc_hd__xor2_1
X_1027_ _1054_/A _1054_/B _1041_/B _1026_/X VGND VGND VPWR VPWR _1085_/B sky130_fd_sc_hd__o211ai_4
XFILLER_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1714_ _1714_/A VGND VGND VPWR VPWR _1838_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1576_ _1576_/A VGND VGND VPWR VPWR _1763_/D sky130_fd_sc_hd__clkbuf_1
X_1645_ _1645_/A VGND VGND VPWR VPWR _1776_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_58_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1430_ _1155_/A _1428_/Y _1429_/X VGND VGND VPWR VPWR _1431_/B sky130_fd_sc_hd__o21ai_2
XFILLER_48_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1292_ _1446_/A _1279_/B _1271_/B VGND VGND VPWR VPWR _1294_/B sky130_fd_sc_hd__a21o_1
X_1361_ _1361_/A _1381_/A _1361_/C VGND VGND VPWR VPWR _1361_/X sky130_fd_sc_hd__or3_1
XFILLER_63_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1559_ _1559_/A VGND VGND VPWR VPWR _1666_/A sky130_fd_sc_hd__clkinv_2
X_1628_ _1628_/A _1628_/B VGND VGND VPWR VPWR _1628_/Y sky130_fd_sc_hd__nand2_1
XTAP_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0930_ _0910_/Y _0920_/X _1287_/A VGND VGND VPWR VPWR _0931_/A sky130_fd_sc_hd__mux2_1
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1413_ _1447_/B _1413_/B VGND VGND VPWR VPWR _1413_/X sky130_fd_sc_hd__xor2_1
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1344_ _1344_/A _1344_/B VGND VGND VPWR VPWR _1357_/A sky130_fd_sc_hd__nor2_1
X_1275_ _0972_/B _1220_/B _1273_/X _1274_/X VGND VGND VPWR VPWR _1448_/A sky130_fd_sc_hd__a211o_1
XFILLER_36_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1060_ _1060_/A _1060_/B VGND VGND VPWR VPWR _1060_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_18_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0913_ _0937_/A VGND VGND VPWR VPWR _1020_/A sky130_fd_sc_hd__inv_2
XFILLER_64_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1327_ _1327_/A VGND VGND VPWR VPWR _1420_/A sky130_fd_sc_hd__clkbuf_2
X_1258_ _1313_/A _1258_/B VGND VGND VPWR VPWR _1260_/B sky130_fd_sc_hd__nand2_1
X_1189_ _1212_/B _1188_/X _1173_/X VGND VGND VPWR VPWR _1190_/C sky130_fd_sc_hd__a21bo_1
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1043_ _1069_/A _1069_/C _1043_/C _1043_/D VGND VGND VPWR VPWR _1047_/C sky130_fd_sc_hd__or4_1
XFILLER_53_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1112_ _1112_/A VGND VGND VPWR VPWR _1220_/B sky130_fd_sc_hd__buf_2
XFILLER_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1592_ _1613_/B VGND VGND VPWR VPWR _1624_/B sky130_fd_sc_hd__clkbuf_2
X_1661_ _1661_/A VGND VGND VPWR VPWR _1781_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1730_ _1730_/A VGND VGND VPWR VPWR _1845_/D sky130_fd_sc_hd__clkbuf_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1026_ _1205_/B _1026_/B VGND VGND VPWR VPWR _1026_/X sky130_fd_sc_hd__or2_1
XFILLER_53_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1713_ _1785_/Q _1554_/A input4/X VGND VGND VPWR VPWR _1714_/A sky130_fd_sc_hd__mux2_1
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1575_ _1762_/Q _1575_/B VGND VGND VPWR VPWR _1576_/A sky130_fd_sc_hd__and2_1
X_1644_ _1647_/A _1644_/B VGND VGND VPWR VPWR _1645_/A sky130_fd_sc_hd__and2_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_0 input2/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1009_ _1221_/B _1026_/B VGND VGND VPWR VPWR _1054_/A sky130_fd_sc_hd__xnor2_2
XFILLER_34_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1360_ _1360_/A _1360_/B _1360_/C VGND VGND VPWR VPWR _1361_/C sky130_fd_sc_hd__and3_1
X_1291_ _1291_/A _1291_/B VGND VGND VPWR VPWR _1446_/B sky130_fd_sc_hd__nor2_1
XFILLER_23_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1627_ _1627_/A _1627_/B VGND VGND VPWR VPWR _1628_/B sky130_fd_sc_hd__xnor2_1
X_1558_ _1558_/A VGND VGND VPWR VPWR _1667_/B sky130_fd_sc_hd__clkbuf_2
XTAP_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1489_ _1495_/B VGND VGND VPWR VPWR _1504_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1343_ _1180_/A _1341_/B _1342_/Y _1339_/X VGND VGND VPWR VPWR _1344_/B sky130_fd_sc_hd__o2bb2a_1
X_1412_ _1411_/Y _1371_/B _1329_/B VGND VGND VPWR VPWR _1413_/B sky130_fd_sc_hd__o21ai_1
XFILLER_5_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1274_ _0972_/B _1220_/B _1206_/A VGND VGND VPWR VPWR _1274_/X sky130_fd_sc_hd__o21a_1
XFILLER_36_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0989_ _0979_/B _0981_/Y _1008_/S VGND VGND VPWR VPWR _0991_/B sky130_fd_sc_hd__mux2_1
XFILLER_59_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0912_ _1392_/A _0937_/A _0910_/B VGND VGND VPWR VPWR _0919_/A sky130_fd_sc_hd__or3b_1
XFILLER_18_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1326_ _1392_/A _1422_/B VGND VGND VPWR VPWR _1329_/A sky130_fd_sc_hd__nand2_1
XFILLER_64_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1257_ _1257_/A _1257_/B _1257_/C VGND VGND VPWR VPWR _1258_/B sky130_fd_sc_hd__or3_1
X_1188_ _1277_/C _1315_/A VGND VGND VPWR VPWR _1188_/X sky130_fd_sc_hd__or2b_1
XFILLER_17_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1042_ _1085_/A _1041_/B _1041_/C VGND VGND VPWR VPWR _1043_/D sky130_fd_sc_hd__a21oi_1
X_1111_ _1290_/B _1106_/X _1110_/X _1249_/B VGND VGND VPWR VPWR _1111_/X sky130_fd_sc_hd__o22a_1
XFILLER_46_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1309_ _1310_/A _1310_/B VGND VGND VPWR VPWR _1360_/B sky130_fd_sc_hd__nand2_1
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1591_ _1582_/X _1584_/X _1585_/Y _1583_/X VGND VGND VPWR VPWR _1613_/B sky130_fd_sc_hd__o22a_1
X_1660_ _1675_/A _1660_/B VGND VGND VPWR VPWR _1661_/A sky130_fd_sc_hd__and2_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1025_ _1221_/B VGND VGND VPWR VPWR _1205_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_53_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1789_ _1789_/D _1551_/Y VGND VGND VPWR VPWR _1789_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_55_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1712_ _1712_/A VGND VGND VPWR VPWR _1837_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1643_ _1776_/Q _1814_/Q _1650_/S VGND VGND VPWR VPWR _1644_/B sky130_fd_sc_hd__mux2_1
XFILLER_39_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1574_ _1574_/A VGND VGND VPWR VPWR _1762_/D sky130_fd_sc_hd__clkbuf_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1008_ _1005_/Y _1007_/Y _1008_/S VGND VGND VPWR VPWR _1026_/B sky130_fd_sc_hd__mux2_2
XFILLER_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1290_ _1290_/A _1290_/B VGND VGND VPWR VPWR _1291_/B sky130_fd_sc_hd__nor2_1
XFILLER_36_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1626_ _1545_/A _1620_/B _1625_/X VGND VGND VPWR VPWR _1627_/B sky130_fd_sc_hd__o21a_1
X_1557_ _1668_/B _1668_/C VGND VGND VPWR VPWR _1558_/A sky130_fd_sc_hd__and2_1
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1488_ _1774_/Q _1778_/Q _1835_/Q VGND VGND VPWR VPWR _1495_/B sky130_fd_sc_hd__mux2_1
XFILLER_52_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1342_ _1342_/A VGND VGND VPWR VPWR _1342_/Y sky130_fd_sc_hd__clkinv_2
X_1273_ _1273_/A _1276_/A _1281_/A _1273_/D VGND VGND VPWR VPWR _1273_/X sky130_fd_sc_hd__and4_1
X_1411_ _1420_/A _1411_/B VGND VGND VPWR VPWR _1411_/Y sky130_fd_sc_hd__nor2_1
XFILLER_51_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0988_ _0988_/A _0988_/B VGND VGND VPWR VPWR _1008_/S sky130_fd_sc_hd__nor2_2
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1609_ _1607_/X _1609_/B _1609_/C VGND VGND VPWR VPWR _1609_/X sky130_fd_sc_hd__and3b_1
XFILLER_47_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_0911_ _1828_/Q VGND VGND VPWR VPWR _0937_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1256_ _1257_/A _1257_/B _1257_/C VGND VGND VPWR VPWR _1313_/A sky130_fd_sc_hd__o21ai_1
X_1325_ _1193_/X _1287_/X _1321_/X _1324_/Y _1217_/X VGND VGND VPWR VPWR _1791_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_64_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1187_ _1272_/B _1273_/A _1315_/A VGND VGND VPWR VPWR _1212_/B sky130_fd_sc_hd__a21o_1
XFILLER_33_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1110_ _1107_/X _1109_/Y _1149_/S VGND VGND VPWR VPWR _1110_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1041_ _1085_/A _1041_/B _1041_/C VGND VGND VPWR VPWR _1043_/C sky130_fd_sc_hd__and3_1
XFILLER_46_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1308_ _1338_/A _1308_/B VGND VGND VPWR VPWR _1310_/B sky130_fd_sc_hd__xnor2_1
X_1239_ _1276_/A _1209_/B _1206_/B VGND VGND VPWR VPWR _1240_/B sky130_fd_sc_hd__a21oi_1
XFILLER_29_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1590_ _1534_/A _1588_/X _1589_/Y VGND VGND VPWR VPWR _1766_/D sky130_fd_sc_hd__o21a_1
X_1024_ _1112_/A _1024_/B VGND VGND VPWR VPWR _1041_/B sky130_fd_sc_hd__or2_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1788_ _1788_/D _1551_/Y VGND VGND VPWR VPWR _1788_/Q sky130_fd_sc_hd__dlxtn_1
X_1857_ _1816_/Q _1857_/D VGND VGND VPWR VPWR _1857_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1711_ _1784_/Q _1532_/B _1711_/S VGND VGND VPWR VPWR _1712_/A sky130_fd_sc_hd__mux2_1
XFILLER_6_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1642_ _1642_/A VGND VGND VPWR VPWR _1775_/D sky130_fd_sc_hd__clkbuf_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1573_ _1761_/Q _1575_/B VGND VGND VPWR VPWR _1574_/A sky130_fd_sc_hd__and2_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1007_ _1007_/A _1007_/B VGND VGND VPWR VPWR _1007_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_34_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1556_ _1556_/A VGND VGND VPWR VPWR _1668_/C sky130_fd_sc_hd__inv_2
X_1625_ _1771_/Q _1624_/B _1619_/X VGND VGND VPWR VPWR _1625_/X sky130_fd_sc_hd__a21bo_1
XFILLER_39_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1487_ _1777_/Q _1708_/B _1482_/X VGND VGND VPWR VPWR _1498_/C sky130_fd_sc_hd__o21ai_1
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1410_ _1409_/A _1409_/B _1409_/C VGND VGND VPWR VPWR _1410_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1341_ _1339_/X _1341_/B _1341_/C _1342_/A VGND VGND VPWR VPWR _1344_/A sky130_fd_sc_hd__and4b_1
X_1272_ _1277_/B _1272_/B VGND VGND VPWR VPWR _1273_/D sky130_fd_sc_hd__nand2_1
X_0987_ _0985_/A _0947_/Y _0907_/B VGND VGND VPWR VPWR _0988_/B sky130_fd_sc_hd__a21o_1
XFILLER_59_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1539_ _1539_/A VGND VGND VPWR VPWR _1821_/D sky130_fd_sc_hd__clkbuf_1
X_1608_ _1768_/Q _1807_/D _1806_/D _1613_/B VGND VGND VPWR VPWR _1609_/B sky130_fd_sc_hd__a31o_1
XFILLER_63_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_0910_ _1327_/A _0910_/B VGND VGND VPWR VPWR _0910_/Y sky130_fd_sc_hd__nand2_1
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1255_ _1255_/A _1255_/B VGND VGND VPWR VPWR _1257_/C sky130_fd_sc_hd__xnor2_1
X_1186_ _1149_/S _1287_/B _1173_/X _1185_/X VGND VGND VPWR VPWR _1190_/B sky130_fd_sc_hd__a211o_1
X_1324_ _1322_/Y _1323_/X _1193_/A VGND VGND VPWR VPWR _1324_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_32_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1040_ _1054_/A _1054_/B _1026_/X VGND VGND VPWR VPWR _1041_/C sky130_fd_sc_hd__o21a_1
XFILLER_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1307_ _1346_/A _1346_/B VGND VGND VPWR VPWR _1308_/B sky130_fd_sc_hd__xor2_1
XFILLER_37_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1238_ _1238_/A _1238_/B VGND VGND VPWR VPWR _1238_/X sky130_fd_sc_hd__xor2_1
X_1169_ _1690_/A VGND VGND VPWR VPWR _1735_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1023_ _1060_/A _1059_/B _1022_/X VGND VGND VPWR VPWR _1054_/B sky130_fd_sc_hd__a21oi_4
XFILLER_38_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1787_ _1787_/D _1551_/Y VGND VGND VPWR VPWR _1787_/Q sky130_fd_sc_hd__dlxtn_1
X_1856_ _1816_/Q _1856_/D VGND VGND VPWR VPWR _1856_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1710_ _1710_/A VGND VGND VPWR VPWR _1836_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1641_ _1647_/A _1641_/B VGND VGND VPWR VPWR _1642_/A sky130_fd_sc_hd__and2_1
X_1572_ _1572_/A VGND VGND VPWR VPWR _1761_/D sky130_fd_sc_hd__clkbuf_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1006_ _1350_/B _1006_/B VGND VGND VPWR VPWR _1007_/B sky130_fd_sc_hd__xnor2_1
XFILLER_26_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1839_ _1839_/CLK _1840_/Q VGND VGND VPWR VPWR _1839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1624_ _1772_/Q _1624_/B VGND VGND VPWR VPWR _1627_/A sky130_fd_sc_hd__xor2_1
X_1555_ _1555_/A VGND VGND VPWR VPWR _1555_/X sky130_fd_sc_hd__clkbuf_1
XTAP_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1486_ _1498_/B VGND VGND VPWR VPWR _1505_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_62_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1340_ _1339_/A _1327_/A _1821_/Q _1339_/D VGND VGND VPWR VPWR _1342_/A sky130_fd_sc_hd__a22o_1
X_1271_ _1271_/A _1271_/B VGND VGND VPWR VPWR _1446_/A sky130_fd_sc_hd__nor2_2
XFILLER_36_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_0986_ _1028_/B _1028_/C _1028_/A VGND VGND VPWR VPWR _0988_/A sky130_fd_sc_hd__a21oi_2
X_1538_ _1603_/A _1538_/B VGND VGND VPWR VPWR _1539_/A sky130_fd_sc_hd__and2_1
X_1607_ _1768_/Q _1807_/D _1806_/D _1613_/B VGND VGND VPWR VPWR _1607_/X sky130_fd_sc_hd__o31a_1
X_1469_ _1769_/Q VGND VGND VPWR VPWR _1541_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_63_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1323_ _1426_/C _1323_/B _1446_/B VGND VGND VPWR VPWR _1323_/X sky130_fd_sc_hd__and3_1
XFILLER_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1254_ _1225_/B _1345_/A _1253_/X VGND VGND VPWR VPWR _1255_/B sky130_fd_sc_hd__a21oi_1
X_1185_ _1208_/B _1178_/Y _1210_/A _1184_/X VGND VGND VPWR VPWR _1185_/X sky130_fd_sc_hd__a31o_1
XFILLER_24_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_0969_ _1244_/A _1244_/B _1823_/Q VGND VGND VPWR VPWR _1004_/B sky130_fd_sc_hd__a21o_1
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1306_ _1345_/A _1345_/B _1305_/X VGND VGND VPWR VPWR _1346_/B sky130_fd_sc_hd__o21ai_1
XFILLER_64_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1099_ _1101_/A _1101_/C VGND VGND VPWR VPWR _1100_/C sky130_fd_sc_hd__nor2_1
XFILLER_52_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1237_ _1246_/A _1245_/A VGND VGND VPWR VPWR _1238_/B sky130_fd_sc_hd__nand2_1
X_1168_ _1727_/B VGND VGND VPWR VPWR _1690_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_12_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1022_ _1392_/B _1057_/A _1057_/B VGND VGND VPWR VPWR _1022_/X sky130_fd_sc_hd__and3_1
XFILLER_19_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1855_ _1816_/Q _1855_/D VGND VGND VPWR VPWR _1855_/Q sky130_fd_sc_hd__dfxtp_1
X_1786_ _1786_/D _1551_/Y VGND VGND VPWR VPWR _1786_/Q sky130_fd_sc_hd__dlxtn_1
XFILLER_55_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1571_ _1760_/Q _1575_/B VGND VGND VPWR VPWR _1572_/A sky130_fd_sc_hd__and2_1
X_1640_ _1775_/Q _1813_/Q _1650_/S VGND VGND VPWR VPWR _1641_/B sky130_fd_sc_hd__mux2_1
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_1005_ _1006_/B VGND VGND VPWR VPWR _1005_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1838_ _1839_/CLK _1838_/D VGND VGND VPWR VPWR _1838_/Q sky130_fd_sc_hd__dfxtp_1
X_1769_ _1816_/Q _1769_/D VGND VGND VPWR VPWR _1769_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput6 _1804_/Q VGND VGND VPWR VPWR led_flag sky130_fd_sc_hd__buf_2
XFILLER_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1623_ _1545_/A _1588_/X _1622_/X _1599_/X VGND VGND VPWR VPWR _1771_/D sky130_fd_sc_hd__o211a_1
X_1554_ _1554_/A VGND VGND VPWR VPWR _1555_/A sky130_fd_sc_hd__clkbuf_1
XTAP_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1485_ _1485_/A _1505_/B VGND VGND VPWR VPWR _1485_/Y sky130_fd_sc_hd__nand2_1
.ends

