* NGSPICE file created from PrimitiveCalculator.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

.subckt PrimitiveCalculator VGND VPWR clk led_flag restart rotary_a rotary_b rst select
+ seven_segment_digit seven_segment_out[0] seven_segment_out[1] seven_segment_out[2]
+ seven_segment_out[3] seven_segment_out[4] seven_segment_out[5] seven_segment_out[6]
XFILLER_36_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_13__4 VGND VGND VPWR VPWR _13__4/HI seven_segment_out[6] sky130_fd_sc_hd__conb_1
XFILLER_63_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_08__7 VGND VGND VPWR VPWR seven_segment_out[2] _08__7/LO sky130_fd_sc_hd__conb_1
XFILLER_5_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_10__9 VGND VGND VPWR VPWR seven_segment_out[4] _10__9/LO sky130_fd_sc_hd__conb_1
XFILLER_37_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_05_ _04_/Q _05_/D VGND VGND VPWR VPWR _05_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_04_ clk _04_/D VGND VGND VPWR VPWR _04_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput1 rst VGND VGND VPWR VPWR _03_/B sky130_fd_sc_hd__buf_2
XFILLER_36_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_03_ _05_/Q _03_/B VGND VGND VPWR VPWR _05_/D sky130_fd_sc_hd__nor2_1
XFILLER_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_02_ _04_/Q _03_/B VGND VGND VPWR VPWR _04_/D sky130_fd_sc_hd__nor2_1
XFILLER_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_06__5 VGND VGND VPWR VPWR seven_segment_out[0] _06__5/LO sky130_fd_sc_hd__conb_1
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_09__8 VGND VGND VPWR VPWR seven_segment_out[3] _09__8/LO sky130_fd_sc_hd__conb_1
XFILLER_0_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_12__3 VGND VGND VPWR VPWR _12__3/HI led_flag sky130_fd_sc_hd__conb_1
XFILLER_36_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_07__6 VGND VGND VPWR VPWR seven_segment_out[1] _07__6/LO sky130_fd_sc_hd__conb_1
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput2 _05_/Q VGND VGND VPWR VPWR seven_segment_digit sky130_fd_sc_hd__buf_2
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_11__10 VGND VGND VPWR VPWR seven_segment_out[5] _11__10/LO sky130_fd_sc_hd__conb_1
XFILLER_40_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

