magic
tech sky130A
magscale 1 2
timestamp 1651670678
<< viali >>
rect 25237 37417 25271 37451
rect 23857 37349 23891 37383
rect 25329 37349 25363 37383
rect 25881 37349 25915 37383
rect 25237 37281 25271 37315
rect 27353 37281 27387 37315
rect 28549 37281 28583 37315
rect 3801 37213 3835 37247
rect 14105 37213 14139 37247
rect 23673 37213 23707 37247
rect 25421 37213 25455 37247
rect 26157 37213 26191 37247
rect 26341 37213 26375 37247
rect 28641 37213 28675 37247
rect 30297 37213 30331 37247
rect 30481 37213 30515 37247
rect 34713 37213 34747 37247
rect 25053 37145 25087 37179
rect 26985 37145 27019 37179
rect 27169 37145 27203 37179
rect 28273 37145 28307 37179
rect 28733 37145 28767 37179
rect 3985 37077 4019 37111
rect 14289 37077 14323 37111
rect 26065 37077 26099 37111
rect 28365 37077 28399 37111
rect 30389 37077 30423 37111
rect 34897 37077 34931 37111
rect 25421 36873 25455 36907
rect 28825 36873 28859 36907
rect 29745 36873 29779 36907
rect 24409 36805 24443 36839
rect 25329 36805 25363 36839
rect 26249 36805 26283 36839
rect 24225 36737 24259 36771
rect 24501 36737 24535 36771
rect 26157 36737 26191 36771
rect 26341 36737 26375 36771
rect 27445 36737 27479 36771
rect 28641 36737 28675 36771
rect 28917 36737 28951 36771
rect 29653 36737 29687 36771
rect 29837 36737 29871 36771
rect 30481 36737 30515 36771
rect 25605 36669 25639 36703
rect 27537 36669 27571 36703
rect 28457 36669 28491 36703
rect 30573 36669 30607 36703
rect 24225 36601 24259 36635
rect 24961 36533 24995 36567
rect 27721 36533 27755 36567
rect 30757 36533 30791 36567
rect 23765 36329 23799 36363
rect 24961 36329 24995 36363
rect 26249 36329 26283 36363
rect 29837 36329 29871 36363
rect 30665 36329 30699 36363
rect 30941 36329 30975 36363
rect 31585 36329 31619 36363
rect 25145 36261 25179 36295
rect 30021 36261 30055 36295
rect 26249 36193 26283 36227
rect 28733 36193 28767 36227
rect 28825 36193 28859 36227
rect 31493 36193 31527 36227
rect 32597 36193 32631 36227
rect 23673 36125 23707 36159
rect 26157 36125 26191 36159
rect 26433 36125 26467 36159
rect 29653 36125 29687 36159
rect 29745 36125 29779 36159
rect 30481 36125 30515 36159
rect 31401 36125 31435 36159
rect 31677 36125 31711 36159
rect 32321 36125 32355 36159
rect 32413 36125 32447 36159
rect 24777 36057 24811 36091
rect 24977 35989 25011 36023
rect 26617 35989 26651 36023
rect 28273 35989 28307 36023
rect 28641 35989 28675 36023
rect 31861 35989 31895 36023
rect 32597 35989 32631 36023
rect 24777 35785 24811 35819
rect 26341 35785 26375 35819
rect 27445 35785 27479 35819
rect 29485 35785 29519 35819
rect 29653 35785 29687 35819
rect 32505 35785 32539 35819
rect 25973 35717 26007 35751
rect 27353 35717 27387 35751
rect 28733 35717 28767 35751
rect 29285 35717 29319 35751
rect 23581 35649 23615 35683
rect 23765 35649 23799 35683
rect 24961 35649 24995 35683
rect 25053 35649 25087 35683
rect 25237 35649 25271 35683
rect 25329 35649 25363 35683
rect 26157 35649 26191 35683
rect 26433 35649 26467 35683
rect 28273 35649 28307 35683
rect 28457 35649 28491 35683
rect 31125 35649 31159 35683
rect 31309 35649 31343 35683
rect 31585 35649 31619 35683
rect 32137 35649 32171 35683
rect 32965 35649 32999 35683
rect 33149 35649 33183 35683
rect 27537 35581 27571 35615
rect 28825 35581 28859 35615
rect 31217 35581 31251 35615
rect 32229 35581 32263 35615
rect 23673 35445 23707 35479
rect 26985 35445 27019 35479
rect 29469 35445 29503 35479
rect 30849 35445 30883 35479
rect 31401 35445 31435 35479
rect 32321 35445 32355 35479
rect 33057 35445 33091 35479
rect 24409 35241 24443 35275
rect 27169 35241 27203 35275
rect 28641 35241 28675 35275
rect 29653 35241 29687 35275
rect 31953 35241 31987 35275
rect 25881 35173 25915 35207
rect 27813 35173 27847 35207
rect 27353 35105 27387 35139
rect 30941 35105 30975 35139
rect 20177 35037 20211 35071
rect 20361 35037 20395 35071
rect 20821 35037 20855 35071
rect 21005 35037 21039 35071
rect 23673 35037 23707 35071
rect 23857 35037 23891 35071
rect 24567 35037 24601 35071
rect 24674 35037 24708 35071
rect 24777 35037 24811 35071
rect 24869 35037 24903 35071
rect 25789 35037 25823 35071
rect 26065 35037 26099 35071
rect 26249 35037 26283 35071
rect 26525 35037 26559 35071
rect 27077 35037 27111 35071
rect 27813 35037 27847 35071
rect 28089 35037 28123 35071
rect 28549 35037 28583 35071
rect 28733 35037 28767 35071
rect 29929 35037 29963 35071
rect 31585 35037 31619 35071
rect 31769 35037 31803 35071
rect 29653 34969 29687 35003
rect 29837 34969 29871 35003
rect 30849 34969 30883 35003
rect 20269 34901 20303 34935
rect 20913 34901 20947 34935
rect 23857 34901 23891 34935
rect 27353 34901 27387 34935
rect 27997 34901 28031 34935
rect 30389 34901 30423 34935
rect 30757 34901 30791 34935
rect 19625 34697 19659 34731
rect 21833 34697 21867 34731
rect 26249 34697 26283 34731
rect 30573 34697 30607 34731
rect 31401 34697 31435 34731
rect 24409 34629 24443 34663
rect 28457 34629 28491 34663
rect 28657 34629 28691 34663
rect 30205 34629 30239 34663
rect 30405 34629 30439 34663
rect 19441 34561 19475 34595
rect 19625 34561 19659 34595
rect 20269 34561 20303 34595
rect 21097 34561 21131 34595
rect 21189 34561 21223 34595
rect 22201 34561 22235 34595
rect 24869 34561 24903 34595
rect 26157 34561 26191 34595
rect 26341 34561 26375 34595
rect 26985 34561 27019 34595
rect 27169 34561 27203 34595
rect 27629 34561 27663 34595
rect 27813 34561 27847 34595
rect 29285 34561 29319 34595
rect 29469 34561 29503 34595
rect 31033 34561 31067 34595
rect 31217 34561 31251 34595
rect 32137 34561 32171 34595
rect 37841 34561 37875 34595
rect 20361 34493 20395 34527
rect 22293 34493 22327 34527
rect 22477 34493 22511 34527
rect 23581 34493 23615 34527
rect 25145 34493 25179 34527
rect 27077 34493 27111 34527
rect 32413 34493 32447 34527
rect 20637 34425 20671 34459
rect 27997 34357 28031 34391
rect 28641 34357 28675 34391
rect 28825 34357 28859 34391
rect 29285 34357 29319 34391
rect 30389 34357 30423 34391
rect 32229 34357 32263 34391
rect 32321 34357 32355 34391
rect 38025 34357 38059 34391
rect 19809 34153 19843 34187
rect 21649 34153 21683 34187
rect 28181 34153 28215 34187
rect 28641 34153 28675 34187
rect 29837 34153 29871 34187
rect 30021 34153 30055 34187
rect 31309 34153 31343 34187
rect 19993 34085 20027 34119
rect 26157 34085 26191 34119
rect 32965 34085 32999 34119
rect 20637 34017 20671 34051
rect 23857 34017 23891 34051
rect 25513 34017 25547 34051
rect 26709 34017 26743 34051
rect 28365 34017 28399 34051
rect 29653 34017 29687 34051
rect 33057 34017 33091 34051
rect 19625 33949 19659 33983
rect 19809 33949 19843 33983
rect 20453 33949 20487 33983
rect 20821 33949 20855 33983
rect 21465 33949 21499 33983
rect 23489 33949 23523 33983
rect 23765 33949 23799 33983
rect 24685 33949 24719 33983
rect 24869 33949 24903 33983
rect 25145 33949 25179 33983
rect 25973 33949 26007 33983
rect 26985 33949 27019 33983
rect 28181 33949 28215 33983
rect 28457 33949 28491 33983
rect 29837 33949 29871 33983
rect 30481 33949 30515 33983
rect 30665 33949 30699 33983
rect 31125 33949 31159 33983
rect 31309 33949 31343 33983
rect 31953 33949 31987 33983
rect 32137 33949 32171 33983
rect 32781 33949 32815 33983
rect 32873 33949 32907 33983
rect 21281 33881 21315 33915
rect 29561 33881 29595 33915
rect 32321 33881 32355 33915
rect 20545 33813 20579 33847
rect 20729 33813 20763 33847
rect 30573 33813 30607 33847
rect 31493 33813 31527 33847
rect 24961 33609 24995 33643
rect 26985 33609 27019 33643
rect 30297 33609 30331 33643
rect 20453 33541 20487 33575
rect 24133 33541 24167 33575
rect 31217 33541 31251 33575
rect 19349 33473 19383 33507
rect 19625 33473 19659 33507
rect 20269 33473 20303 33507
rect 20361 33473 20395 33507
rect 20637 33473 20671 33507
rect 20729 33473 20763 33507
rect 22201 33473 22235 33507
rect 23949 33473 23983 33507
rect 24041 33473 24075 33507
rect 24317 33473 24351 33507
rect 24409 33473 24443 33507
rect 24869 33473 24903 33507
rect 25053 33473 25087 33507
rect 25881 33473 25915 33507
rect 27169 33473 27203 33507
rect 27445 33473 27479 33507
rect 28457 33473 28491 33507
rect 28733 33473 28767 33507
rect 29101 33473 29135 33507
rect 29929 33473 29963 33507
rect 30113 33473 30147 33507
rect 30941 33473 30975 33507
rect 31089 33473 31123 33507
rect 31309 33473 31343 33507
rect 31425 33473 31459 33507
rect 32505 33473 32539 33507
rect 33977 33473 34011 33507
rect 22293 33405 22327 33439
rect 22477 33405 22511 33439
rect 25605 33405 25639 33439
rect 27353 33405 27387 33439
rect 28181 33405 28215 33439
rect 32781 33405 32815 33439
rect 33885 33405 33919 33439
rect 19165 33337 19199 33371
rect 28733 33337 28767 33371
rect 34345 33337 34379 33371
rect 19533 33269 19567 33303
rect 20085 33269 20119 33303
rect 21833 33269 21867 33303
rect 23765 33269 23799 33303
rect 31585 33269 31619 33303
rect 20637 33065 20671 33099
rect 23857 33065 23891 33099
rect 25329 33065 25363 33099
rect 25881 33065 25915 33099
rect 28181 33065 28215 33099
rect 30021 33065 30055 33099
rect 30205 33065 30239 33099
rect 33057 33065 33091 33099
rect 17601 32997 17635 33031
rect 21833 32997 21867 33031
rect 24685 32997 24719 33031
rect 26985 32997 27019 33031
rect 31677 32997 31711 33031
rect 20821 32929 20855 32963
rect 21373 32929 21407 32963
rect 23489 32929 23523 32963
rect 26157 32929 26191 32963
rect 26249 32929 26283 32963
rect 29837 32929 29871 32963
rect 31125 32929 31159 32963
rect 33517 32929 33551 32963
rect 33701 32929 33735 32963
rect 34805 32929 34839 32963
rect 1409 32861 1443 32895
rect 16773 32861 16807 32895
rect 17049 32861 17083 32895
rect 17233 32861 17267 32895
rect 18061 32861 18095 32895
rect 20361 32861 20395 32895
rect 21465 32861 21499 32895
rect 22293 32861 22327 32895
rect 22477 32861 22511 32895
rect 23673 32861 23707 32895
rect 24409 32861 24443 32895
rect 24685 32861 24719 32895
rect 25237 32861 25271 32895
rect 25421 32861 25455 32895
rect 26065 32861 26099 32895
rect 26341 32861 26375 32895
rect 26525 32861 26559 32895
rect 27169 32861 27203 32895
rect 27445 32861 27479 32895
rect 28365 32861 28399 32895
rect 28549 32861 28583 32895
rect 28641 32861 28675 32895
rect 30021 32861 30055 32895
rect 31677 32861 31711 32895
rect 31861 32861 31895 32895
rect 32321 32861 32355 32895
rect 32505 32861 32539 32895
rect 32597 32861 32631 32895
rect 32689 32861 32723 32895
rect 32873 32861 32907 32895
rect 33793 32861 33827 32895
rect 33885 32861 33919 32895
rect 33977 32861 34011 32895
rect 34897 32861 34931 32895
rect 17601 32793 17635 32827
rect 29561 32793 29595 32827
rect 30849 32793 30883 32827
rect 1593 32725 1627 32759
rect 18153 32725 18187 32759
rect 22385 32725 22419 32759
rect 27353 32725 27387 32759
rect 35265 32725 35299 32759
rect 16865 32521 16899 32555
rect 18547 32521 18581 32555
rect 19349 32521 19383 32555
rect 21113 32521 21147 32555
rect 23581 32521 23615 32555
rect 25973 32521 26007 32555
rect 29193 32521 29227 32555
rect 33793 32521 33827 32555
rect 18337 32453 18371 32487
rect 20913 32453 20947 32487
rect 24409 32453 24443 32487
rect 27353 32453 27387 32487
rect 30297 32453 30331 32487
rect 30507 32453 30541 32487
rect 33701 32453 33735 32487
rect 15761 32385 15795 32419
rect 17049 32385 17083 32419
rect 17325 32385 17359 32419
rect 17509 32385 17543 32419
rect 19290 32385 19324 32419
rect 22569 32385 22603 32419
rect 22845 32385 22879 32419
rect 23029 32385 23063 32419
rect 23489 32385 23523 32419
rect 23673 32385 23707 32419
rect 24317 32385 24351 32419
rect 24501 32385 24535 32419
rect 25145 32385 25179 32419
rect 26157 32385 26191 32419
rect 26341 32385 26375 32419
rect 26433 32385 26467 32419
rect 27169 32385 27203 32419
rect 27445 32385 27479 32419
rect 28181 32385 28215 32419
rect 28549 32385 28583 32419
rect 30205 32385 30239 32419
rect 30389 32385 30423 32419
rect 31309 32385 31343 32419
rect 31493 32385 31527 32419
rect 32137 32385 32171 32419
rect 32321 32385 32355 32419
rect 32597 32385 32631 32419
rect 15669 32317 15703 32351
rect 17233 32317 17267 32351
rect 19809 32317 19843 32351
rect 24961 32317 24995 32351
rect 30665 32317 30699 32351
rect 31585 32317 31619 32351
rect 32689 32317 32723 32351
rect 33885 32317 33919 32351
rect 16129 32249 16163 32283
rect 17141 32249 17175 32283
rect 21281 32249 21315 32283
rect 22385 32249 22419 32283
rect 18521 32181 18555 32215
rect 18705 32181 18739 32215
rect 19165 32181 19199 32215
rect 19717 32181 19751 32215
rect 21097 32181 21131 32215
rect 25329 32181 25363 32215
rect 26985 32181 27019 32215
rect 30021 32181 30055 32215
rect 31125 32181 31159 32215
rect 33333 32181 33367 32215
rect 15301 31977 15335 32011
rect 16313 31977 16347 32011
rect 16957 31977 16991 32011
rect 20637 31977 20671 32011
rect 23213 31977 23247 32011
rect 24777 31977 24811 32011
rect 26893 31977 26927 32011
rect 33517 31977 33551 32011
rect 18521 31909 18555 31943
rect 24961 31909 24995 31943
rect 25605 31909 25639 31943
rect 28641 31909 28675 31943
rect 15945 31841 15979 31875
rect 17049 31841 17083 31875
rect 18245 31841 18279 31875
rect 18705 31841 18739 31875
rect 19349 31841 19383 31875
rect 21741 31841 21775 31875
rect 22293 31841 22327 31875
rect 23673 31841 23707 31875
rect 26065 31841 26099 31875
rect 29561 31841 29595 31875
rect 34069 31841 34103 31875
rect 15301 31773 15335 31807
rect 15485 31773 15519 31807
rect 16129 31773 16163 31807
rect 16773 31773 16807 31807
rect 16865 31773 16899 31807
rect 19441 31773 19475 31807
rect 20821 31773 20855 31807
rect 21097 31773 21131 31807
rect 21925 31773 21959 31807
rect 26157 31773 26191 31807
rect 26801 31773 26835 31807
rect 28273 31773 28307 31807
rect 28457 31773 28491 31807
rect 29837 31773 29871 31807
rect 31217 31773 31251 31807
rect 31309 31773 31343 31807
rect 31401 31773 31435 31807
rect 31585 31773 31619 31807
rect 32229 31773 32263 31807
rect 32321 31773 32355 31807
rect 32505 31773 32539 31807
rect 32597 31773 32631 31807
rect 33149 31773 33183 31807
rect 33333 31773 33367 31807
rect 33977 31773 34011 31807
rect 34161 31773 34195 31807
rect 34713 31773 34747 31807
rect 34897 31773 34931 31807
rect 17601 31705 17635 31739
rect 23765 31705 23799 31739
rect 24593 31705 24627 31739
rect 27629 31705 27663 31739
rect 27813 31705 27847 31739
rect 17693 31637 17727 31671
rect 19809 31637 19843 31671
rect 21005 31637 21039 31671
rect 22201 31637 22235 31671
rect 23673 31637 23707 31671
rect 24793 31637 24827 31671
rect 26065 31637 26099 31671
rect 30941 31637 30975 31671
rect 32045 31637 32079 31671
rect 34805 31637 34839 31671
rect 15209 31433 15243 31467
rect 16129 31433 16163 31467
rect 16865 31433 16899 31467
rect 18337 31433 18371 31467
rect 18797 31433 18831 31467
rect 19165 31433 19199 31467
rect 21833 31433 21867 31467
rect 24593 31433 24627 31467
rect 29193 31433 29227 31467
rect 33149 31433 33183 31467
rect 17969 31365 18003 31399
rect 18185 31365 18219 31399
rect 21097 31365 21131 31399
rect 27261 31365 27295 31399
rect 15117 31297 15151 31331
rect 15301 31297 15335 31331
rect 15945 31297 15979 31331
rect 17049 31297 17083 31331
rect 17141 31297 17175 31331
rect 17325 31297 17359 31331
rect 18981 31297 19015 31331
rect 19257 31297 19291 31331
rect 20085 31297 20119 31331
rect 20361 31297 20395 31331
rect 21005 31297 21039 31331
rect 21189 31297 21223 31331
rect 22109 31297 22143 31331
rect 23029 31297 23063 31331
rect 23857 31297 23891 31331
rect 24041 31297 24075 31331
rect 24501 31297 24535 31331
rect 25605 31297 25639 31331
rect 25881 31297 25915 31331
rect 26157 31297 26191 31331
rect 26341 31297 26375 31331
rect 26985 31297 27019 31331
rect 27078 31297 27112 31331
rect 27353 31297 27387 31331
rect 27491 31297 27525 31331
rect 28273 31297 28307 31331
rect 28365 31297 28399 31331
rect 28641 31297 28675 31331
rect 29101 31297 29135 31331
rect 29929 31297 29963 31331
rect 30573 31297 30607 31331
rect 30757 31297 30791 31331
rect 30941 31297 30975 31331
rect 31125 31297 31159 31331
rect 32781 31297 32815 31331
rect 33609 31297 33643 31331
rect 33793 31297 33827 31331
rect 34529 31297 34563 31331
rect 35541 31297 35575 31331
rect 15761 31229 15795 31263
rect 20177 31229 20211 31263
rect 22017 31229 22051 31263
rect 22201 31229 22235 31263
rect 22293 31229 22327 31263
rect 22937 31229 22971 31263
rect 25973 31229 26007 31263
rect 29745 31229 29779 31263
rect 30849 31229 30883 31263
rect 32689 31229 32723 31263
rect 34621 31229 34655 31263
rect 34897 31229 34931 31263
rect 35449 31229 35483 31263
rect 17233 31161 17267 31195
rect 20545 31161 20579 31195
rect 28549 31161 28583 31195
rect 33609 31161 33643 31195
rect 35909 31161 35943 31195
rect 18153 31093 18187 31127
rect 20085 31093 20119 31127
rect 23305 31093 23339 31127
rect 23949 31093 23983 31127
rect 27629 31093 27663 31127
rect 28089 31093 28123 31127
rect 30113 31093 30147 31127
rect 31309 31093 31343 31127
rect 15209 30889 15243 30923
rect 16405 30889 16439 30923
rect 20729 30889 20763 30923
rect 21281 30889 21315 30923
rect 29745 30889 29779 30923
rect 30665 30889 30699 30923
rect 31125 30889 31159 30923
rect 31493 30889 31527 30923
rect 31585 30889 31619 30923
rect 32505 30889 32539 30923
rect 32689 30889 32723 30923
rect 33425 30889 33459 30923
rect 18153 30821 18187 30855
rect 19257 30821 19291 30855
rect 23489 30821 23523 30855
rect 25237 30821 25271 30855
rect 31401 30821 31435 30855
rect 23213 30753 23247 30787
rect 28273 30753 28307 30787
rect 36001 30753 36035 30787
rect 15485 30685 15519 30719
rect 15577 30685 15611 30719
rect 15669 30685 15703 30719
rect 15853 30685 15887 30719
rect 16589 30685 16623 30719
rect 16865 30685 16899 30719
rect 17049 30685 17083 30719
rect 17785 30685 17819 30719
rect 17969 30685 18003 30719
rect 18153 30685 18187 30719
rect 18521 30685 18555 30719
rect 19441 30685 19475 30719
rect 19717 30685 19751 30719
rect 20453 30685 20487 30719
rect 20545 30685 20579 30719
rect 21465 30685 21499 30719
rect 21741 30685 21775 30719
rect 22201 30685 22235 30719
rect 22385 30685 22419 30719
rect 23121 30685 23155 30719
rect 26065 30685 26099 30719
rect 26249 30685 26283 30719
rect 26893 30685 26927 30719
rect 26985 30685 27019 30719
rect 27169 30685 27203 30719
rect 27261 30685 27295 30719
rect 28181 30685 28215 30719
rect 28733 30685 28767 30719
rect 30297 30685 30331 30719
rect 31677 30685 31711 30719
rect 31861 30685 31895 30719
rect 32321 30685 32355 30719
rect 32505 30685 32539 30719
rect 33425 30685 33459 30719
rect 33609 30685 33643 30719
rect 35081 30685 35115 30719
rect 35265 30685 35299 30719
rect 35909 30685 35943 30719
rect 16681 30617 16715 30651
rect 16773 30617 16807 30651
rect 24961 30617 24995 30651
rect 29653 30617 29687 30651
rect 30481 30617 30515 30651
rect 19625 30549 19659 30583
rect 21649 30549 21683 30583
rect 22293 30549 22327 30583
rect 25421 30549 25455 30583
rect 26157 30549 26191 30583
rect 26709 30549 26743 30583
rect 28917 30549 28951 30583
rect 35173 30549 35207 30583
rect 36277 30549 36311 30583
rect 18521 30345 18555 30379
rect 18981 30345 19015 30379
rect 22201 30345 22235 30379
rect 22871 30345 22905 30379
rect 34897 30345 34931 30379
rect 15761 30277 15795 30311
rect 20821 30277 20855 30311
rect 22661 30277 22695 30311
rect 23765 30277 23799 30311
rect 27721 30277 27755 30311
rect 32321 30277 32355 30311
rect 33977 30277 34011 30311
rect 15577 30209 15611 30243
rect 15853 30209 15887 30243
rect 15945 30209 15979 30243
rect 16681 30209 16715 30243
rect 17049 30209 17083 30243
rect 17417 30209 17451 30243
rect 18245 30209 18279 30243
rect 19257 30209 19291 30243
rect 19441 30209 19475 30243
rect 20085 30209 20119 30243
rect 20729 30209 20763 30243
rect 21833 30209 21867 30243
rect 22017 30209 22051 30243
rect 23581 30209 23615 30243
rect 24501 30209 24535 30243
rect 25237 30209 25271 30243
rect 25881 30209 25915 30243
rect 27629 30209 27663 30243
rect 27813 30209 27847 30243
rect 27951 30209 27985 30243
rect 28733 30209 28767 30243
rect 31401 30209 31435 30243
rect 32137 30209 32171 30243
rect 32413 30209 32447 30243
rect 32873 30209 32907 30243
rect 33057 30209 33091 30243
rect 34161 30209 34195 30243
rect 34897 30209 34931 30243
rect 36277 30209 36311 30243
rect 37473 30209 37507 30243
rect 17785 30141 17819 30175
rect 19165 30141 19199 30175
rect 19349 30141 19383 30175
rect 20269 30141 20303 30175
rect 24317 30141 24351 30175
rect 25973 30141 26007 30175
rect 28089 30141 28123 30175
rect 30021 30141 30055 30175
rect 30297 30141 30331 30175
rect 31585 30141 31619 30175
rect 34437 30141 34471 30175
rect 35173 30141 35207 30175
rect 36185 30141 36219 30175
rect 37381 30141 37415 30175
rect 16129 30073 16163 30107
rect 25421 30073 25455 30107
rect 27445 30073 27479 30107
rect 34345 30073 34379 30107
rect 34989 30073 35023 30107
rect 37841 30073 37875 30107
rect 22845 30005 22879 30039
rect 23029 30005 23063 30039
rect 24685 30005 24719 30039
rect 28917 30005 28951 30039
rect 32137 30005 32171 30039
rect 32873 30005 32907 30039
rect 36553 30005 36587 30039
rect 15945 29801 15979 29835
rect 18061 29801 18095 29835
rect 18337 29801 18371 29835
rect 19993 29801 20027 29835
rect 21281 29801 21315 29835
rect 22937 29801 22971 29835
rect 24593 29801 24627 29835
rect 26341 29801 26375 29835
rect 36093 29801 36127 29835
rect 25697 29733 25731 29767
rect 26525 29733 26559 29767
rect 33701 29733 33735 29767
rect 16681 29665 16715 29699
rect 24501 29665 24535 29699
rect 24685 29665 24719 29699
rect 25421 29665 25455 29699
rect 27813 29665 27847 29699
rect 30205 29665 30239 29699
rect 31861 29665 31895 29699
rect 32137 29665 32171 29699
rect 33241 29665 33275 29699
rect 15577 29597 15611 29631
rect 16405 29597 16439 29631
rect 17969 29597 18003 29631
rect 18153 29597 18187 29631
rect 21097 29597 21131 29631
rect 22661 29597 22695 29631
rect 23397 29597 23431 29631
rect 23581 29597 23615 29631
rect 24409 29597 24443 29631
rect 25329 29597 25363 29631
rect 28641 29597 28675 29631
rect 31033 29597 31067 29631
rect 33333 29597 33367 29631
rect 34713 29597 34747 29631
rect 34897 29597 34931 29631
rect 35357 29597 35391 29631
rect 35541 29597 35575 29631
rect 36093 29597 36127 29631
rect 36369 29597 36403 29631
rect 15761 29529 15795 29563
rect 19809 29529 19843 29563
rect 22385 29529 22419 29563
rect 22569 29529 22603 29563
rect 26157 29529 26191 29563
rect 30021 29529 30055 29563
rect 30849 29529 30883 29563
rect 36277 29529 36311 29563
rect 20009 29461 20043 29495
rect 20177 29461 20211 29495
rect 22753 29461 22787 29495
rect 23673 29461 23707 29495
rect 26357 29461 26391 29495
rect 34805 29461 34839 29495
rect 35449 29461 35483 29495
rect 17417 29257 17451 29291
rect 17785 29257 17819 29291
rect 23029 29257 23063 29291
rect 27445 29257 27479 29291
rect 28089 29257 28123 29291
rect 28749 29257 28783 29291
rect 31309 29257 31343 29291
rect 32337 29257 32371 29291
rect 32505 29257 32539 29291
rect 33241 29257 33275 29291
rect 37933 29257 37967 29291
rect 16773 29189 16807 29223
rect 16957 29189 16991 29223
rect 28549 29189 28583 29223
rect 29653 29189 29687 29223
rect 32137 29189 32171 29223
rect 36461 29189 36495 29223
rect 15945 29121 15979 29155
rect 16129 29121 16163 29155
rect 17601 29121 17635 29155
rect 17877 29121 17911 29155
rect 18337 29121 18371 29155
rect 18521 29121 18555 29155
rect 19533 29121 19567 29155
rect 19717 29121 19751 29155
rect 19901 29121 19935 29155
rect 20269 29121 20303 29155
rect 20729 29121 20763 29155
rect 22293 29121 22327 29155
rect 22937 29121 22971 29155
rect 23121 29121 23155 29155
rect 23857 29121 23891 29155
rect 23949 29121 23983 29155
rect 24092 29121 24126 29155
rect 24235 29121 24269 29155
rect 24869 29121 24903 29155
rect 25053 29121 25087 29155
rect 25145 29121 25179 29155
rect 26065 29121 26099 29155
rect 29469 29121 29503 29155
rect 29745 29121 29779 29155
rect 29837 29121 29871 29155
rect 30481 29121 30515 29155
rect 30665 29121 30699 29155
rect 31217 29121 31251 29155
rect 32965 29121 32999 29155
rect 33885 29121 33919 29155
rect 34713 29121 34747 29155
rect 35725 29121 35759 29155
rect 36645 29121 36679 29155
rect 36737 29121 36771 29155
rect 26249 29053 26283 29087
rect 27813 29053 27847 29087
rect 27905 29053 27939 29087
rect 33241 29053 33275 29087
rect 33977 29053 34011 29087
rect 34805 29053 34839 29087
rect 35541 29053 35575 29087
rect 37289 29053 37323 29087
rect 37657 29053 37691 29087
rect 37749 29053 37783 29087
rect 16037 28985 16071 29019
rect 22477 28985 22511 29019
rect 28917 28985 28951 29019
rect 30573 28985 30607 29019
rect 34253 28985 34287 29019
rect 35081 28985 35115 29019
rect 36737 28985 36771 29019
rect 18429 28917 18463 28951
rect 19533 28917 19567 28951
rect 20821 28917 20855 28951
rect 23673 28917 23707 28951
rect 24685 28917 24719 28951
rect 28733 28917 28767 28951
rect 30021 28917 30055 28951
rect 32321 28917 32355 28951
rect 33057 28917 33091 28951
rect 34805 28917 34839 28951
rect 35909 28917 35943 28951
rect 15485 28713 15519 28747
rect 16957 28713 16991 28747
rect 18521 28713 18555 28747
rect 19809 28713 19843 28747
rect 21925 28713 21959 28747
rect 23857 28713 23891 28747
rect 24961 28713 24995 28747
rect 27721 28713 27755 28747
rect 31953 28713 31987 28747
rect 34897 28713 34931 28747
rect 36829 28713 36863 28747
rect 37933 28713 37967 28747
rect 18705 28645 18739 28679
rect 21005 28645 21039 28679
rect 17601 28577 17635 28611
rect 20063 28577 20097 28611
rect 20168 28577 20202 28611
rect 28457 28577 28491 28611
rect 34069 28577 34103 28611
rect 34805 28577 34839 28611
rect 34989 28577 35023 28611
rect 15669 28509 15703 28543
rect 16313 28509 16347 28543
rect 17325 28509 17359 28543
rect 19967 28509 20001 28543
rect 20262 28509 20296 28543
rect 20821 28509 20855 28543
rect 21005 28509 21039 28543
rect 21833 28509 21867 28543
rect 22017 28509 22051 28543
rect 22845 28509 22879 28543
rect 23029 28509 23063 28543
rect 24869 28509 24903 28543
rect 26065 28509 26099 28543
rect 26341 28509 26375 28543
rect 27189 28509 27223 28543
rect 27537 28509 27571 28543
rect 28181 28509 28215 28543
rect 30849 28509 30883 28543
rect 31033 28509 31067 28543
rect 32137 28509 32171 28543
rect 32229 28509 32263 28543
rect 32689 28509 32723 28543
rect 32873 28509 32907 28543
rect 33333 28509 33367 28543
rect 33517 28509 33551 28543
rect 33977 28509 34011 28543
rect 34161 28509 34195 28543
rect 34713 28509 34747 28543
rect 35817 28509 35851 28543
rect 37013 28509 37047 28543
rect 37197 28509 37231 28543
rect 37289 28509 37323 28543
rect 16129 28441 16163 28475
rect 16497 28441 16531 28475
rect 17417 28441 17451 28475
rect 18337 28441 18371 28475
rect 21373 28441 21407 28475
rect 23489 28441 23523 28475
rect 23673 28441 23707 28475
rect 26433 28441 26467 28475
rect 27353 28441 27387 28475
rect 27445 28441 27479 28475
rect 30021 28441 30055 28475
rect 31953 28441 31987 28475
rect 33425 28441 33459 28475
rect 36001 28441 36035 28475
rect 37749 28441 37783 28475
rect 37949 28441 37983 28475
rect 18547 28373 18581 28407
rect 30113 28373 30147 28407
rect 30941 28373 30975 28407
rect 32781 28373 32815 28407
rect 36185 28373 36219 28407
rect 38117 28373 38151 28407
rect 17325 28169 17359 28203
rect 18521 28169 18555 28203
rect 23397 28169 23431 28203
rect 28457 28169 28491 28203
rect 30113 28169 30147 28203
rect 31401 28169 31435 28203
rect 34437 28169 34471 28203
rect 37657 28169 37691 28203
rect 16957 28101 16991 28135
rect 17173 28101 17207 28135
rect 18889 28101 18923 28135
rect 20821 28101 20855 28135
rect 31125 28101 31159 28135
rect 32413 28101 32447 28135
rect 33885 28101 33919 28135
rect 15117 28033 15151 28067
rect 17877 28033 17911 28067
rect 18705 28033 18739 28067
rect 18981 28033 19015 28067
rect 19809 28033 19843 28067
rect 19901 28033 19935 28067
rect 20637 28033 20671 28067
rect 20729 28033 20763 28067
rect 21005 28033 21039 28067
rect 21097 28033 21131 28067
rect 21833 28033 21867 28067
rect 22569 28033 22603 28067
rect 23213 28033 23247 28067
rect 24041 28033 24075 28067
rect 24777 28033 24811 28067
rect 24961 28033 24995 28067
rect 25789 28033 25823 28067
rect 25973 28033 26007 28067
rect 27445 28033 27479 28067
rect 28365 28033 28399 28067
rect 29101 28033 29135 28067
rect 29285 28033 29319 28067
rect 29377 28033 29411 28067
rect 29837 28033 29871 28067
rect 30849 28033 30883 28067
rect 31033 28033 31067 28067
rect 31217 28033 31251 28067
rect 32137 28033 32171 28067
rect 32229 28033 32263 28067
rect 32505 28033 32539 28067
rect 32597 28033 32631 28067
rect 33701 28033 33735 28067
rect 34345 28033 34379 28067
rect 34529 28033 34563 28067
rect 34989 28033 35023 28067
rect 35173 28033 35207 28067
rect 35909 28033 35943 28067
rect 36093 28033 36127 28067
rect 36553 28033 36587 28067
rect 36737 28033 36771 28067
rect 37473 28033 37507 28067
rect 37749 28033 37783 28067
rect 14841 27965 14875 27999
rect 19441 27965 19475 27999
rect 19625 27965 19659 27999
rect 19717 27965 19751 27999
rect 30113 27965 30147 27999
rect 20453 27897 20487 27931
rect 22753 27897 22787 27931
rect 27629 27897 27663 27931
rect 32137 27897 32171 27931
rect 36001 27897 36035 27931
rect 15853 27829 15887 27863
rect 17141 27829 17175 27863
rect 17969 27829 18003 27863
rect 21925 27829 21959 27863
rect 24133 27829 24167 27863
rect 25881 27829 25915 27863
rect 29929 27829 29963 27863
rect 34989 27829 35023 27863
rect 36645 27829 36679 27863
rect 37473 27829 37507 27863
rect 16957 27625 16991 27659
rect 18153 27625 18187 27659
rect 19441 27625 19475 27659
rect 19993 27625 20027 27659
rect 21189 27625 21223 27659
rect 25881 27625 25915 27659
rect 27629 27625 27663 27659
rect 28325 27625 28359 27659
rect 16405 27557 16439 27591
rect 34713 27557 34747 27591
rect 36645 27557 36679 27591
rect 23029 27489 23063 27523
rect 29837 27489 29871 27523
rect 32137 27489 32171 27523
rect 32413 27489 32447 27523
rect 34161 27489 34195 27523
rect 35541 27489 35575 27523
rect 36185 27489 36219 27523
rect 14473 27421 14507 27455
rect 14749 27421 14783 27455
rect 16221 27421 16255 27455
rect 16957 27421 16991 27455
rect 17233 27421 17267 27455
rect 17785 27421 17819 27455
rect 18061 27421 18095 27455
rect 20177 27421 20211 27455
rect 20453 27421 20487 27455
rect 21833 27421 21867 27455
rect 22017 27421 22051 27455
rect 23213 27421 23247 27455
rect 24869 27421 24903 27455
rect 26525 27421 26559 27455
rect 27169 27421 27203 27455
rect 27353 27421 27387 27455
rect 29653 27421 29687 27455
rect 30297 27421 30331 27455
rect 30481 27421 30515 27455
rect 30941 27421 30975 27455
rect 32229 27421 32263 27455
rect 32321 27421 32355 27455
rect 33642 27421 33676 27455
rect 34069 27421 34103 27455
rect 34713 27421 34747 27455
rect 35449 27421 35483 27455
rect 35633 27421 35667 27455
rect 36277 27421 36311 27455
rect 37105 27421 37139 27455
rect 37289 27421 37323 27455
rect 37749 27421 37783 27455
rect 37933 27421 37967 27455
rect 19349 27353 19383 27387
rect 21097 27353 21131 27387
rect 25789 27353 25823 27387
rect 27721 27353 27755 27387
rect 28181 27353 28215 27387
rect 37197 27353 37231 27387
rect 15485 27285 15519 27319
rect 17141 27285 17175 27319
rect 18337 27285 18371 27319
rect 20361 27285 20395 27319
rect 22201 27285 22235 27319
rect 23397 27285 23431 27319
rect 25145 27285 25179 27319
rect 26617 27285 26651 27319
rect 28381 27285 28415 27319
rect 28549 27285 28583 27319
rect 30389 27285 30423 27319
rect 31033 27285 31067 27319
rect 31953 27285 31987 27319
rect 33517 27285 33551 27319
rect 33701 27285 33735 27319
rect 37841 27285 37875 27319
rect 15393 27081 15427 27115
rect 20361 27081 20395 27115
rect 25053 27081 25087 27115
rect 25973 27081 26007 27115
rect 28825 27081 28859 27115
rect 33517 27081 33551 27115
rect 33793 27081 33827 27115
rect 36553 27081 36587 27115
rect 18061 27013 18095 27047
rect 19625 27013 19659 27047
rect 21097 27013 21131 27047
rect 21281 27013 21315 27047
rect 23673 27013 23707 27047
rect 28457 27013 28491 27047
rect 29929 27013 29963 27047
rect 32505 27013 32539 27047
rect 33425 27013 33459 27047
rect 14657 26945 14691 26979
rect 15945 26945 15979 26979
rect 16129 26945 16163 26979
rect 16773 26945 16807 26979
rect 19441 26945 19475 26979
rect 19717 26945 19751 26979
rect 20177 26945 20211 26979
rect 20453 26945 20487 26979
rect 22385 26945 22419 26979
rect 22661 26945 22695 26979
rect 23489 26945 23523 26979
rect 24133 26945 24167 26979
rect 24225 26945 24259 26979
rect 24961 26945 24995 26979
rect 25145 26945 25179 26979
rect 25605 26945 25639 26979
rect 25789 26945 25823 26979
rect 28273 26945 28307 26979
rect 28549 26945 28583 26979
rect 28687 26945 28721 26979
rect 29653 26945 29687 26979
rect 29837 26945 29871 26979
rect 30021 26945 30055 26979
rect 31150 26945 31184 26979
rect 32321 26945 32355 26979
rect 32413 26945 32447 26979
rect 32689 26945 32723 26979
rect 33149 26945 33183 26979
rect 34621 26945 34655 26979
rect 34713 26945 34747 26979
rect 34805 26945 34839 26979
rect 34989 26945 35023 26979
rect 35725 26945 35759 26979
rect 35909 26945 35943 26979
rect 36461 26945 36495 26979
rect 36645 26945 36679 26979
rect 37473 26945 37507 26979
rect 14381 26877 14415 26911
rect 16865 26877 16899 26911
rect 22753 26877 22787 26911
rect 22937 26877 22971 26911
rect 26985 26877 27019 26911
rect 27261 26877 27295 26911
rect 30665 26877 30699 26911
rect 30941 26877 30975 26911
rect 31033 26877 31067 26911
rect 33634 26877 33668 26911
rect 35633 26877 35667 26911
rect 35817 26877 35851 26911
rect 37381 26877 37415 26911
rect 17693 26809 17727 26843
rect 20177 26809 20211 26843
rect 32137 26809 32171 26843
rect 15945 26741 15979 26775
rect 16865 26741 16899 26775
rect 17141 26741 17175 26775
rect 18061 26741 18095 26775
rect 18245 26741 18279 26775
rect 19257 26741 19291 26775
rect 30205 26741 30239 26775
rect 31309 26741 31343 26775
rect 34345 26741 34379 26775
rect 35449 26741 35483 26775
rect 37749 26741 37783 26775
rect 16773 26537 16807 26571
rect 17785 26537 17819 26571
rect 25053 26537 25087 26571
rect 26709 26537 26743 26571
rect 27261 26537 27295 26571
rect 35909 26537 35943 26571
rect 36185 26537 36219 26571
rect 18337 26469 18371 26503
rect 19717 26469 19751 26503
rect 26065 26469 26099 26503
rect 26617 26469 26651 26503
rect 28549 26469 28583 26503
rect 33057 26469 33091 26503
rect 14197 26401 14231 26435
rect 18061 26401 18095 26435
rect 21465 26401 21499 26435
rect 21833 26401 21867 26435
rect 23305 26401 23339 26435
rect 26801 26401 26835 26435
rect 30757 26401 30791 26435
rect 32045 26401 32079 26435
rect 33977 26401 34011 26435
rect 34713 26401 34747 26435
rect 14473 26333 14507 26367
rect 15301 26333 15335 26367
rect 15761 26333 15795 26367
rect 16037 26333 16071 26367
rect 17693 26333 17727 26367
rect 18153 26333 18187 26367
rect 19901 26333 19935 26367
rect 19993 26333 20027 26367
rect 20177 26333 20211 26367
rect 20269 26333 20303 26367
rect 21557 26333 21591 26367
rect 21925 26333 21959 26367
rect 23213 26333 23247 26367
rect 24961 26333 24995 26367
rect 25881 26333 25915 26367
rect 26525 26333 26559 26367
rect 27445 26333 27479 26367
rect 27537 26333 27571 26367
rect 27721 26333 27755 26367
rect 27813 26333 27847 26367
rect 29561 26333 29595 26367
rect 29745 26333 29779 26367
rect 30481 26333 30515 26367
rect 30573 26333 30607 26367
rect 30849 26333 30883 26367
rect 32505 26333 32539 26367
rect 32781 26333 32815 26367
rect 32873 26333 32907 26367
rect 34897 26333 34931 26367
rect 34989 26333 35023 26367
rect 35173 26333 35207 26367
rect 35265 26333 35299 26367
rect 35725 26333 35759 26367
rect 37289 26333 37323 26367
rect 37749 26333 37783 26367
rect 21281 26265 21315 26299
rect 23857 26265 23891 26299
rect 28365 26265 28399 26299
rect 29653 26265 29687 26299
rect 30297 26265 30331 26299
rect 31861 26265 31895 26299
rect 32689 26265 32723 26299
rect 33793 26265 33827 26299
rect 38117 26265 38151 26299
rect 21741 26197 21775 26231
rect 13185 25993 13219 26027
rect 14473 25993 14507 26027
rect 16129 25993 16163 26027
rect 17693 25993 17727 26027
rect 18337 25993 18371 26027
rect 22569 25993 22603 26027
rect 30573 25993 30607 26027
rect 33701 25993 33735 26027
rect 35357 25993 35391 26027
rect 18245 25925 18279 25959
rect 24133 25925 24167 25959
rect 27445 25925 27479 25959
rect 27629 25925 27663 25959
rect 29377 25925 29411 25959
rect 29593 25925 29627 25959
rect 32597 25925 32631 25959
rect 33333 25925 33367 25959
rect 33517 25925 33551 25959
rect 35265 25925 35299 25959
rect 36093 25925 36127 25959
rect 13369 25857 13403 25891
rect 14013 25857 14047 25891
rect 14657 25857 14691 25891
rect 15393 25857 15427 25891
rect 16957 25857 16991 25891
rect 18889 25857 18923 25891
rect 19901 25857 19935 25891
rect 20269 25857 20303 25891
rect 20729 25857 20763 25891
rect 20913 25857 20947 25891
rect 22385 25857 22419 25891
rect 23121 25857 23155 25891
rect 24041 25857 24075 25891
rect 24225 25857 24259 25891
rect 24869 25857 24903 25891
rect 25881 25857 25915 25891
rect 26157 25857 26191 25891
rect 26341 25857 26375 25891
rect 27721 25857 27755 25891
rect 28549 25857 28583 25891
rect 30389 25857 30423 25891
rect 30665 25857 30699 25891
rect 31125 25857 31159 25891
rect 31309 25857 31343 25891
rect 32321 25857 32355 25891
rect 32505 25857 32539 25891
rect 32689 25857 32723 25891
rect 33609 25857 33643 25891
rect 34345 25857 34379 25891
rect 35909 25857 35943 25891
rect 36185 25857 36219 25891
rect 37473 25857 37507 25891
rect 15117 25789 15151 25823
rect 16681 25789 16715 25823
rect 19717 25789 19751 25823
rect 20821 25789 20855 25823
rect 24961 25789 24995 25823
rect 25053 25789 25087 25823
rect 25145 25789 25179 25823
rect 28733 25789 28767 25823
rect 28825 25789 28859 25823
rect 30205 25789 30239 25823
rect 37565 25789 37599 25823
rect 13829 25721 13863 25755
rect 20177 25721 20211 25755
rect 23305 25721 23339 25755
rect 25973 25721 26007 25755
rect 26065 25721 26099 25755
rect 27445 25721 27479 25755
rect 29745 25721 29779 25755
rect 19073 25653 19107 25687
rect 24685 25653 24719 25687
rect 25697 25653 25731 25687
rect 28365 25653 28399 25687
rect 29561 25653 29595 25687
rect 31217 25653 31251 25687
rect 32873 25653 32907 25687
rect 33885 25653 33919 25687
rect 34529 25653 34563 25687
rect 35909 25653 35943 25687
rect 37749 25653 37783 25687
rect 13369 25449 13403 25483
rect 14105 25449 14139 25483
rect 15117 25449 15151 25483
rect 15761 25449 15795 25483
rect 17417 25449 17451 25483
rect 20637 25449 20671 25483
rect 22109 25449 22143 25483
rect 30757 25449 30791 25483
rect 34713 25449 34747 25483
rect 36001 25449 36035 25483
rect 21189 25381 21223 25415
rect 22753 25381 22787 25415
rect 25697 25381 25731 25415
rect 29837 25381 29871 25415
rect 16405 25313 16439 25347
rect 22845 25313 22879 25347
rect 23673 25313 23707 25347
rect 23857 25313 23891 25347
rect 33333 25313 33367 25347
rect 35357 25313 35391 25347
rect 37565 25313 37599 25347
rect 13553 25245 13587 25279
rect 14289 25245 14323 25279
rect 15301 25245 15335 25279
rect 15945 25245 15979 25279
rect 16681 25245 16715 25279
rect 18613 25245 18647 25279
rect 19625 25245 19659 25279
rect 19901 25245 19935 25279
rect 21097 25245 21131 25279
rect 22477 25245 22511 25279
rect 22569 25245 22603 25279
rect 23581 25245 23615 25279
rect 24409 25245 24443 25279
rect 24685 25245 24719 25279
rect 25973 25245 26007 25279
rect 26893 25245 26927 25279
rect 27077 25245 27111 25279
rect 28181 25245 28215 25279
rect 28273 25245 28307 25279
rect 28457 25245 28491 25279
rect 28549 25245 28583 25279
rect 30113 25245 30147 25279
rect 31585 25245 31619 25279
rect 32505 25245 32539 25279
rect 32689 25245 32723 25279
rect 33609 25245 33643 25279
rect 34838 25245 34872 25279
rect 35265 25245 35299 25279
rect 37473 25245 37507 25279
rect 25697 25177 25731 25211
rect 29837 25177 29871 25211
rect 30573 25177 30607 25211
rect 35817 25177 35851 25211
rect 18429 25109 18463 25143
rect 22391 25109 22425 25143
rect 23857 25109 23891 25143
rect 25881 25109 25915 25143
rect 26985 25109 27019 25143
rect 27997 25109 28031 25143
rect 30021 25109 30055 25143
rect 30773 25109 30807 25143
rect 30941 25109 30975 25143
rect 31401 25109 31435 25143
rect 32597 25109 32631 25143
rect 34897 25109 34931 25143
rect 36017 25109 36051 25143
rect 36185 25109 36219 25143
rect 37841 25109 37875 25143
rect 14565 24905 14599 24939
rect 24593 24905 24627 24939
rect 26433 24905 26467 24939
rect 32873 24905 32907 24939
rect 34069 24905 34103 24939
rect 37289 24905 37323 24939
rect 13369 24837 13403 24871
rect 13569 24837 13603 24871
rect 14197 24837 14231 24871
rect 14397 24837 14431 24871
rect 15025 24837 15059 24871
rect 15225 24837 15259 24871
rect 25421 24837 25455 24871
rect 34989 24837 35023 24871
rect 35909 24837 35943 24871
rect 16129 24769 16163 24803
rect 17141 24769 17175 24803
rect 18613 24769 18647 24803
rect 19993 24769 20027 24803
rect 20453 24769 20487 24803
rect 20545 24769 20579 24803
rect 21097 24769 21131 24803
rect 21281 24769 21315 24803
rect 21833 24769 21867 24803
rect 22109 24769 22143 24803
rect 23397 24769 23431 24803
rect 24409 24769 24443 24803
rect 25605 24769 25639 24803
rect 25697 24769 25731 24803
rect 26157 24769 26191 24803
rect 26985 24769 27019 24803
rect 27169 24769 27203 24803
rect 28089 24769 28123 24803
rect 28917 24769 28951 24803
rect 30573 24769 30607 24803
rect 32137 24769 32171 24803
rect 32321 24769 32355 24803
rect 32781 24769 32815 24803
rect 32965 24769 32999 24803
rect 33701 24769 33735 24803
rect 34186 24769 34220 24803
rect 34823 24769 34857 24803
rect 35173 24769 35207 24803
rect 36093 24769 36127 24803
rect 37473 24769 37507 24803
rect 37657 24769 37691 24803
rect 37749 24769 37783 24803
rect 16865 24701 16899 24735
rect 18337 24701 18371 24735
rect 23673 24701 23707 24735
rect 24225 24701 24259 24735
rect 26433 24701 26467 24735
rect 30389 24701 30423 24735
rect 30757 24701 30791 24735
rect 31217 24701 31251 24735
rect 33977 24701 34011 24735
rect 13737 24633 13771 24667
rect 15393 24633 15427 24667
rect 15945 24633 15979 24667
rect 17877 24633 17911 24667
rect 19809 24633 19843 24667
rect 23489 24633 23523 24667
rect 29285 24633 29319 24667
rect 31125 24633 31159 24667
rect 32229 24633 32263 24667
rect 34345 24633 34379 24667
rect 13553 24565 13587 24599
rect 14381 24565 14415 24599
rect 15209 24565 15243 24599
rect 19349 24565 19383 24599
rect 21189 24565 21223 24599
rect 22845 24565 22879 24599
rect 23581 24565 23615 24599
rect 25421 24565 25455 24599
rect 26249 24565 26283 24599
rect 27353 24565 27387 24599
rect 36277 24565 36311 24599
rect 14289 24361 14323 24395
rect 15117 24361 15151 24395
rect 15945 24361 15979 24395
rect 16129 24361 16163 24395
rect 16773 24361 16807 24395
rect 19809 24361 19843 24395
rect 27537 24361 27571 24395
rect 30481 24361 30515 24395
rect 36737 24361 36771 24395
rect 14473 24293 14507 24327
rect 15301 24293 15335 24327
rect 16957 24293 16991 24327
rect 22017 24293 22051 24327
rect 11529 24225 11563 24259
rect 11989 24225 12023 24259
rect 12541 24225 12575 24259
rect 19441 24225 19475 24259
rect 23305 24225 23339 24259
rect 24593 24225 24627 24259
rect 32505 24225 32539 24259
rect 32965 24225 32999 24259
rect 36369 24225 36403 24259
rect 37289 24225 37323 24259
rect 11621 24157 11655 24191
rect 12633 24157 12667 24191
rect 17509 24157 17543 24191
rect 17693 24157 17727 24191
rect 18521 24157 18555 24191
rect 19625 24157 19659 24191
rect 20361 24157 20395 24191
rect 20545 24157 20579 24191
rect 21005 24157 21039 24191
rect 21281 24157 21315 24191
rect 23213 24157 23247 24191
rect 24501 24157 24535 24191
rect 24685 24157 24719 24191
rect 25145 24157 25179 24191
rect 25329 24157 25363 24191
rect 25789 24157 25823 24191
rect 26801 24157 26835 24191
rect 27077 24157 27111 24191
rect 27537 24157 27571 24191
rect 27721 24157 27755 24191
rect 28733 24157 28767 24191
rect 28917 24157 28951 24191
rect 29561 24157 29595 24191
rect 29745 24157 29779 24191
rect 30389 24157 30423 24191
rect 31217 24157 31251 24191
rect 31401 24157 31435 24191
rect 32229 24157 32263 24191
rect 32321 24157 32355 24191
rect 33241 24157 33275 24191
rect 34713 24157 34747 24191
rect 34897 24157 34931 24191
rect 35357 24157 35391 24191
rect 35541 24157 35575 24191
rect 36553 24157 36587 24191
rect 37381 24157 37415 24191
rect 14105 24089 14139 24123
rect 14310 24089 14344 24123
rect 14933 24089 14967 24123
rect 15761 24089 15795 24123
rect 16589 24089 16623 24123
rect 16789 24089 16823 24123
rect 20453 24089 20487 24123
rect 25881 24089 25915 24123
rect 26985 24089 27019 24123
rect 29929 24089 29963 24123
rect 13001 24021 13035 24055
rect 15133 24021 15167 24055
rect 15961 24021 15995 24055
rect 17877 24021 17911 24055
rect 18337 24021 18371 24055
rect 23581 24021 23615 24055
rect 25237 24021 25271 24055
rect 26617 24021 26651 24055
rect 28825 24021 28859 24055
rect 31309 24021 31343 24055
rect 32505 24021 32539 24055
rect 34805 24021 34839 24055
rect 35541 24021 35575 24055
rect 37749 24021 37783 24055
rect 11897 23817 11931 23851
rect 14289 23817 14323 23851
rect 15777 23817 15811 23851
rect 15945 23817 15979 23851
rect 17969 23817 18003 23851
rect 21189 23817 21223 23851
rect 22109 23817 22143 23851
rect 22753 23817 22787 23851
rect 24409 23817 24443 23851
rect 28917 23817 28951 23851
rect 29101 23817 29135 23851
rect 32505 23817 32539 23851
rect 34897 23817 34931 23851
rect 35817 23817 35851 23851
rect 36461 23817 36495 23851
rect 8585 23749 8619 23783
rect 12265 23749 12299 23783
rect 15577 23749 15611 23783
rect 16865 23749 16899 23783
rect 29653 23749 29687 23783
rect 29837 23749 29871 23783
rect 36277 23749 36311 23783
rect 8401 23681 8435 23715
rect 9229 23681 9263 23715
rect 10149 23681 10183 23715
rect 12081 23681 12115 23715
rect 12357 23681 12391 23715
rect 12817 23681 12851 23715
rect 13001 23681 13035 23715
rect 13461 23681 13495 23715
rect 13645 23681 13679 23715
rect 14473 23681 14507 23715
rect 15117 23681 15151 23715
rect 16681 23681 16715 23715
rect 17785 23681 17819 23715
rect 19165 23681 19199 23715
rect 19993 23681 20027 23715
rect 21097 23681 21131 23715
rect 21281 23681 21315 23715
rect 21925 23681 21959 23715
rect 22109 23681 22143 23715
rect 22569 23681 22603 23715
rect 22753 23681 22787 23715
rect 23397 23681 23431 23715
rect 24225 23681 24259 23715
rect 24409 23681 24443 23715
rect 25421 23681 25455 23715
rect 25605 23681 25639 23715
rect 25697 23681 25731 23715
rect 25881 23681 25915 23715
rect 27261 23681 27295 23715
rect 27445 23681 27479 23715
rect 27905 23681 27939 23715
rect 28089 23681 28123 23715
rect 28733 23681 28767 23715
rect 28825 23681 28859 23715
rect 32413 23681 32447 23715
rect 32597 23681 32631 23715
rect 33057 23681 33091 23715
rect 33241 23681 33275 23715
rect 34529 23681 34563 23715
rect 35357 23681 35391 23715
rect 36553 23681 36587 23715
rect 37473 23681 37507 23715
rect 9321 23613 9355 23647
rect 17601 23613 17635 23647
rect 18981 23613 19015 23647
rect 19809 23613 19843 23647
rect 23305 23613 23339 23647
rect 30665 23613 30699 23647
rect 30941 23613 30975 23647
rect 34621 23613 34655 23647
rect 37565 23613 37599 23647
rect 9597 23545 9631 23579
rect 14933 23545 14967 23579
rect 20177 23545 20211 23579
rect 23765 23545 23799 23579
rect 25513 23545 25547 23579
rect 28549 23545 28583 23579
rect 10241 23477 10275 23511
rect 12817 23477 12851 23511
rect 13553 23477 13587 23511
rect 15761 23477 15795 23511
rect 17049 23477 17083 23511
rect 19349 23477 19383 23511
rect 25237 23477 25271 23511
rect 27353 23477 27387 23511
rect 27997 23477 28031 23511
rect 33149 23477 33183 23511
rect 35449 23477 35483 23511
rect 36277 23477 36311 23511
rect 37841 23477 37875 23511
rect 8401 23273 8435 23307
rect 9505 23273 9539 23307
rect 11621 23273 11655 23307
rect 26065 23273 26099 23307
rect 26801 23273 26835 23307
rect 28549 23273 28583 23307
rect 31493 23273 31527 23307
rect 31861 23273 31895 23307
rect 35909 23273 35943 23307
rect 36737 23273 36771 23307
rect 37105 23273 37139 23307
rect 37657 23273 37691 23307
rect 17785 23205 17819 23239
rect 24777 23205 24811 23239
rect 27721 23205 27755 23239
rect 30849 23205 30883 23239
rect 9229 23137 9263 23171
rect 11161 23137 11195 23171
rect 19625 23137 19659 23171
rect 20453 23137 20487 23171
rect 22017 23137 22051 23171
rect 25513 23137 25547 23171
rect 28457 23137 28491 23171
rect 29745 23137 29779 23171
rect 30389 23137 30423 23171
rect 31585 23137 31619 23171
rect 7021 23069 7055 23103
rect 9137 23069 9171 23103
rect 10241 23069 10275 23103
rect 10333 23069 10367 23103
rect 10425 23069 10459 23103
rect 10609 23069 10643 23103
rect 11253 23069 11287 23103
rect 12725 23069 12759 23103
rect 12817 23069 12851 23103
rect 12909 23069 12943 23103
rect 13093 23069 13127 23103
rect 14105 23069 14139 23103
rect 16773 23069 16807 23103
rect 17049 23069 17083 23103
rect 17601 23069 17635 23103
rect 18705 23069 18739 23103
rect 19257 23069 19291 23103
rect 19441 23069 19475 23103
rect 20729 23069 20763 23103
rect 21557 23069 21591 23103
rect 22293 23069 22327 23103
rect 23581 23069 23615 23103
rect 24777 23069 24811 23103
rect 24961 23069 24995 23103
rect 25421 23069 25455 23103
rect 25605 23069 25639 23103
rect 26341 23069 26375 23103
rect 26801 23069 26835 23103
rect 26985 23069 27019 23103
rect 27629 23069 27663 23103
rect 27813 23069 27847 23103
rect 28273 23069 28307 23103
rect 28549 23069 28583 23103
rect 29653 23069 29687 23103
rect 29837 23069 29871 23103
rect 30481 23069 30515 23103
rect 31493 23069 31527 23103
rect 32781 23069 32815 23103
rect 33701 23069 33735 23103
rect 34897 23069 34931 23103
rect 36645 23069 36679 23103
rect 37565 23069 37599 23103
rect 7288 23001 7322 23035
rect 9965 23001 9999 23035
rect 12449 23001 12483 23035
rect 14350 23001 14384 23035
rect 16589 23001 16623 23035
rect 23765 23001 23799 23035
rect 26065 23001 26099 23035
rect 32965 23001 32999 23035
rect 35081 23001 35115 23035
rect 35725 23001 35759 23035
rect 15485 22933 15519 22967
rect 16957 22933 16991 22967
rect 18521 22933 18555 22967
rect 23029 22933 23063 22967
rect 26249 22933 26283 22967
rect 28733 22933 28767 22967
rect 33149 22933 33183 22967
rect 33793 22933 33827 22967
rect 35265 22933 35299 22967
rect 35925 22933 35959 22967
rect 36093 22933 36127 22967
rect 9597 22729 9631 22763
rect 10609 22729 10643 22763
rect 12357 22729 12391 22763
rect 13093 22729 13127 22763
rect 17601 22729 17635 22763
rect 22661 22729 22695 22763
rect 34621 22729 34655 22763
rect 14289 22661 14323 22695
rect 14841 22661 14875 22695
rect 16681 22661 16715 22695
rect 27353 22661 27387 22695
rect 32229 22661 32263 22695
rect 33609 22661 33643 22695
rect 33825 22661 33859 22695
rect 34437 22661 34471 22695
rect 8769 22593 8803 22627
rect 8953 22593 8987 22627
rect 9045 22593 9079 22627
rect 9781 22593 9815 22627
rect 10057 22593 10091 22627
rect 10517 22593 10551 22627
rect 10701 22593 10735 22627
rect 12173 22593 12207 22627
rect 12817 22593 12851 22627
rect 12909 22593 12943 22627
rect 14105 22593 14139 22627
rect 15577 22593 15611 22627
rect 16865 22593 16899 22627
rect 17785 22593 17819 22627
rect 18429 22593 18463 22627
rect 19073 22593 19107 22627
rect 19257 22593 19291 22627
rect 20269 22593 20303 22627
rect 20545 22593 20579 22627
rect 22753 22593 22787 22627
rect 23489 22593 23523 22627
rect 24501 22593 24535 22627
rect 24593 22593 24627 22627
rect 24777 22593 24811 22627
rect 24869 22593 24903 22627
rect 25697 22593 25731 22627
rect 25789 22593 25823 22627
rect 26985 22593 27019 22627
rect 27078 22593 27112 22627
rect 27261 22593 27295 22627
rect 27491 22593 27525 22627
rect 28365 22593 28399 22627
rect 28549 22593 28583 22627
rect 29193 22593 29227 22627
rect 29377 22593 29411 22627
rect 29837 22593 29871 22627
rect 30021 22593 30055 22627
rect 30573 22593 30607 22627
rect 30757 22593 30791 22627
rect 31217 22593 31251 22627
rect 31309 22593 31343 22627
rect 32137 22593 32171 22627
rect 32321 22593 32355 22627
rect 32965 22593 32999 22627
rect 34713 22593 34747 22627
rect 35357 22593 35391 22627
rect 35449 22593 35483 22627
rect 36093 22593 36127 22627
rect 36277 22593 36311 22627
rect 8861 22525 8895 22559
rect 11989 22525 12023 22559
rect 13093 22525 13127 22559
rect 15025 22525 15059 22559
rect 16957 22525 16991 22559
rect 17049 22525 17083 22559
rect 23581 22525 23615 22559
rect 23857 22525 23891 22559
rect 31493 22525 31527 22559
rect 32781 22525 32815 22559
rect 35633 22525 35667 22559
rect 21281 22457 21315 22491
rect 22385 22457 22419 22491
rect 30573 22457 30607 22491
rect 36461 22457 36495 22491
rect 8585 22389 8619 22423
rect 9965 22389 9999 22423
rect 15577 22389 15611 22423
rect 18245 22389 18279 22423
rect 19441 22389 19475 22423
rect 22017 22389 22051 22423
rect 22293 22389 22327 22423
rect 22477 22389 22511 22423
rect 24317 22389 24351 22423
rect 27629 22389 27663 22423
rect 28733 22389 28767 22423
rect 29285 22389 29319 22423
rect 29929 22389 29963 22423
rect 31401 22389 31435 22423
rect 33149 22389 33183 22423
rect 33793 22389 33827 22423
rect 33977 22389 34011 22423
rect 34437 22389 34471 22423
rect 35541 22389 35575 22423
rect 36277 22389 36311 22423
rect 14841 22185 14875 22219
rect 20729 22185 20763 22219
rect 21649 22185 21683 22219
rect 22661 22185 22695 22219
rect 23029 22185 23063 22219
rect 23673 22185 23707 22219
rect 26249 22185 26283 22219
rect 30573 22185 30607 22219
rect 33149 22185 33183 22219
rect 35541 22185 35575 22219
rect 11161 22117 11195 22151
rect 15485 22117 15519 22151
rect 26985 22117 27019 22151
rect 33517 22117 33551 22151
rect 34805 22117 34839 22151
rect 9505 22049 9539 22083
rect 9965 22049 9999 22083
rect 16405 22049 16439 22083
rect 23121 22049 23155 22083
rect 23857 22049 23891 22083
rect 24961 22049 24995 22083
rect 25145 22049 25179 22083
rect 27169 22049 27203 22083
rect 28089 22049 28123 22083
rect 28273 22049 28307 22083
rect 28365 22049 28399 22083
rect 33609 22049 33643 22083
rect 34989 22049 35023 22083
rect 1409 21981 1443 22015
rect 9597 21981 9631 22015
rect 11877 21981 11911 22015
rect 11970 21981 12004 22015
rect 12102 21981 12136 22015
rect 12265 21981 12299 22015
rect 13553 21981 13587 22015
rect 14197 21981 14231 22015
rect 14381 21981 14415 22015
rect 15025 21981 15059 22015
rect 15485 21981 15519 22015
rect 15669 21981 15703 22015
rect 16129 21981 16163 22015
rect 17417 21981 17451 22015
rect 17785 21981 17819 22015
rect 18705 21981 18739 22015
rect 19257 21981 19291 22015
rect 19441 21981 19475 22015
rect 20269 21981 20303 22015
rect 20913 21981 20947 22015
rect 22845 21981 22879 22015
rect 23581 21981 23615 22015
rect 24409 21981 24443 22015
rect 24869 21981 24903 22015
rect 25237 21981 25271 22015
rect 26157 21981 26191 22015
rect 26893 21981 26927 22015
rect 28181 21981 28215 22015
rect 29561 21981 29595 22015
rect 29745 21981 29779 22015
rect 30205 21981 30239 22015
rect 31217 21981 31251 22015
rect 31401 21981 31435 22015
rect 32413 21981 32447 22015
rect 33333 21981 33367 22015
rect 34713 21981 34747 22015
rect 35449 21981 35483 22015
rect 35633 21981 35667 22015
rect 37381 21981 37415 22015
rect 37749 21981 37783 22015
rect 10977 21913 11011 21947
rect 17601 21913 17635 21947
rect 17693 21913 17727 21947
rect 19625 21913 19659 21947
rect 21465 21913 21499 21947
rect 21681 21913 21715 21947
rect 29653 21913 29687 21947
rect 1593 21845 1627 21879
rect 11621 21845 11655 21879
rect 13369 21845 13403 21879
rect 14381 21845 14415 21879
rect 17969 21845 18003 21879
rect 18521 21845 18555 21879
rect 20085 21845 20119 21879
rect 21833 21845 21867 21879
rect 23857 21845 23891 21879
rect 24501 21845 24535 21879
rect 27169 21845 27203 21879
rect 27905 21845 27939 21879
rect 30573 21845 30607 21879
rect 30757 21845 30791 21879
rect 31309 21845 31343 21879
rect 32505 21845 32539 21879
rect 34713 21845 34747 21879
rect 38117 21845 38151 21879
rect 8677 21641 8711 21675
rect 10609 21641 10643 21675
rect 14381 21641 14415 21675
rect 18153 21641 18187 21675
rect 20085 21641 20119 21675
rect 22753 21641 22787 21675
rect 28917 21641 28951 21675
rect 29653 21641 29687 21675
rect 34069 21641 34103 21675
rect 37841 21641 37875 21675
rect 9321 21573 9355 21607
rect 15393 21573 15427 21607
rect 25789 21573 25823 21607
rect 33701 21573 33735 21607
rect 34529 21573 34563 21607
rect 34713 21573 34747 21607
rect 7564 21505 7598 21539
rect 9689 21505 9723 21539
rect 10517 21505 10551 21539
rect 12173 21505 12207 21539
rect 12265 21505 12299 21539
rect 12449 21505 12483 21539
rect 13001 21505 13035 21539
rect 13268 21505 13302 21539
rect 15301 21505 15335 21539
rect 15945 21505 15979 21539
rect 16129 21505 16163 21539
rect 17141 21505 17175 21539
rect 17436 21505 17470 21539
rect 18613 21505 18647 21539
rect 18889 21505 18923 21539
rect 20269 21505 20303 21539
rect 21005 21505 21039 21539
rect 22569 21505 22603 21539
rect 22845 21505 22879 21539
rect 23305 21505 23339 21539
rect 23489 21505 23523 21539
rect 24133 21505 24167 21539
rect 24317 21505 24351 21539
rect 24961 21505 24995 21539
rect 25053 21505 25087 21539
rect 25237 21505 25271 21539
rect 25329 21505 25363 21539
rect 25973 21505 26007 21539
rect 26065 21505 26099 21539
rect 26249 21505 26283 21539
rect 26341 21505 26375 21539
rect 27445 21505 27479 21539
rect 28733 21505 28767 21539
rect 29009 21505 29043 21539
rect 29469 21505 29503 21539
rect 29745 21505 29779 21539
rect 30849 21505 30883 21539
rect 31033 21505 31067 21539
rect 31125 21505 31159 21539
rect 32137 21505 32171 21539
rect 32321 21505 32355 21539
rect 33885 21505 33919 21539
rect 35633 21505 35667 21539
rect 35909 21505 35943 21539
rect 36093 21505 36127 21539
rect 36369 21505 36403 21539
rect 37473 21505 37507 21539
rect 7297 21437 7331 21471
rect 9781 21437 9815 21471
rect 37565 21437 37599 21471
rect 12357 21369 12391 21403
rect 36185 21369 36219 21403
rect 9965 21301 9999 21335
rect 11989 21301 12023 21335
rect 15945 21301 15979 21335
rect 19625 21301 19659 21335
rect 20821 21301 20855 21335
rect 22385 21301 22419 21335
rect 23673 21301 23707 21335
rect 24133 21301 24167 21335
rect 24777 21301 24811 21335
rect 27721 21301 27755 21335
rect 27905 21301 27939 21335
rect 28549 21301 28583 21335
rect 29469 21301 29503 21335
rect 30665 21301 30699 21335
rect 32137 21301 32171 21335
rect 34897 21301 34931 21335
rect 10149 21097 10183 21131
rect 12817 21097 12851 21131
rect 13461 21097 13495 21131
rect 16681 21097 16715 21131
rect 19257 21097 19291 21131
rect 30021 21097 30055 21131
rect 33333 21097 33367 21131
rect 37013 21097 37047 21131
rect 37657 21097 37691 21131
rect 9505 21029 9539 21063
rect 16313 21029 16347 21063
rect 30573 21029 30607 21063
rect 34897 21029 34931 21063
rect 37565 21029 37599 21063
rect 8401 20961 8435 20995
rect 9689 20961 9723 20995
rect 11437 20961 11471 20995
rect 17693 20961 17727 20995
rect 21833 20961 21867 20995
rect 24777 20961 24811 20995
rect 25053 20961 25087 20995
rect 26893 20961 26927 20995
rect 27353 20961 27387 20995
rect 29653 20961 29687 20995
rect 30757 20961 30791 20995
rect 30849 20961 30883 20995
rect 31033 20961 31067 20995
rect 31585 20961 31619 20995
rect 34989 20961 35023 20995
rect 36737 20961 36771 20995
rect 37749 20961 37783 20995
rect 8125 20893 8159 20927
rect 8217 20893 8251 20927
rect 9413 20893 9447 20927
rect 10425 20893 10459 20927
rect 10517 20893 10551 20927
rect 10609 20893 10643 20927
rect 10793 20893 10827 20927
rect 11704 20893 11738 20927
rect 14473 20893 14507 20927
rect 14729 20893 14763 20927
rect 17969 20893 18003 20927
rect 19441 20893 19475 20927
rect 19901 20893 19935 20927
rect 20177 20893 20211 20927
rect 22109 20893 22143 20927
rect 23351 20893 23385 20927
rect 23486 20890 23520 20924
rect 23581 20893 23615 20927
rect 23765 20893 23799 20927
rect 26249 20893 26283 20927
rect 27261 20893 27295 20927
rect 28365 20893 28399 20927
rect 28825 20893 28859 20927
rect 29009 20893 29043 20927
rect 29745 20893 29779 20927
rect 30941 20893 30975 20927
rect 31769 20893 31803 20927
rect 32413 20893 32447 20927
rect 33241 20893 33275 20927
rect 33333 20893 33367 20927
rect 34713 20893 34747 20927
rect 34805 20893 34839 20927
rect 35633 20893 35667 20927
rect 35725 20893 35759 20927
rect 35909 20893 35943 20927
rect 36001 20893 36035 20927
rect 36645 20893 36679 20927
rect 37473 20893 37507 20927
rect 13369 20825 13403 20859
rect 28089 20825 28123 20859
rect 28273 20825 28307 20859
rect 31953 20825 31987 20859
rect 32597 20825 32631 20859
rect 8401 20757 8435 20791
rect 9689 20757 9723 20791
rect 15853 20757 15887 20791
rect 16681 20757 16715 20791
rect 16865 20757 16899 20791
rect 18705 20757 18739 20791
rect 20913 20757 20947 20791
rect 23121 20757 23155 20791
rect 26341 20757 26375 20791
rect 27537 20757 27571 20791
rect 28187 20757 28221 20791
rect 28917 20757 28951 20791
rect 32781 20757 32815 20791
rect 33609 20757 33643 20791
rect 35449 20757 35483 20791
rect 9965 20553 9999 20587
rect 13185 20553 13219 20587
rect 14841 20553 14875 20587
rect 15301 20553 15335 20587
rect 17325 20553 17359 20587
rect 19257 20553 19291 20587
rect 21833 20553 21867 20587
rect 22937 20553 22971 20587
rect 25897 20553 25931 20587
rect 30205 20553 30239 20587
rect 33149 20553 33183 20587
rect 35541 20553 35575 20587
rect 17233 20485 17267 20519
rect 18429 20485 18463 20519
rect 18889 20485 18923 20519
rect 19089 20485 19123 20519
rect 24961 20485 24995 20519
rect 25697 20485 25731 20519
rect 27353 20485 27387 20519
rect 30113 20485 30147 20519
rect 32689 20485 32723 20519
rect 34989 20485 35023 20519
rect 36369 20485 36403 20519
rect 8677 20417 8711 20451
rect 10149 20417 10183 20451
rect 10333 20417 10367 20451
rect 10425 20417 10459 20451
rect 11897 20417 11931 20451
rect 13369 20417 13403 20451
rect 14105 20417 14139 20451
rect 14289 20417 14323 20451
rect 14381 20417 14415 20451
rect 15209 20417 15243 20451
rect 18061 20417 18095 20451
rect 18245 20417 18279 20451
rect 19993 20417 20027 20451
rect 20269 20417 20303 20451
rect 22017 20417 22051 20451
rect 22109 20417 22143 20451
rect 22293 20417 22327 20451
rect 22477 20417 22511 20451
rect 23121 20417 23155 20451
rect 23949 20417 23983 20451
rect 24225 20417 24259 20451
rect 24409 20417 24443 20451
rect 27077 20417 27111 20451
rect 27170 20417 27204 20451
rect 27445 20417 27479 20451
rect 27583 20417 27617 20451
rect 29009 20417 29043 20451
rect 31217 20417 31251 20451
rect 31401 20417 31435 20451
rect 32232 20417 32266 20451
rect 32505 20417 32539 20451
rect 33517 20417 33551 20451
rect 34253 20417 34287 20451
rect 34437 20417 34471 20451
rect 35725 20417 35759 20451
rect 36185 20417 36219 20451
rect 7573 20349 7607 20383
rect 8769 20349 8803 20383
rect 8861 20349 8895 20383
rect 8953 20349 8987 20383
rect 12173 20349 12207 20383
rect 13645 20349 13679 20383
rect 15485 20349 15519 20383
rect 17509 20349 17543 20383
rect 28733 20349 28767 20383
rect 33609 20349 33643 20383
rect 35449 20349 35483 20383
rect 7941 20281 7975 20315
rect 8493 20281 8527 20315
rect 13553 20281 13587 20315
rect 14105 20281 14139 20315
rect 22201 20281 22235 20315
rect 24041 20281 24075 20315
rect 24133 20281 24167 20315
rect 34989 20281 35023 20315
rect 36553 20281 36587 20315
rect 8033 20213 8067 20247
rect 16865 20213 16899 20247
rect 19073 20213 19107 20247
rect 21005 20213 21039 20247
rect 23765 20213 23799 20247
rect 25053 20213 25087 20247
rect 25881 20213 25915 20247
rect 26065 20213 26099 20247
rect 27721 20213 27755 20247
rect 31585 20213 31619 20247
rect 32597 20213 32631 20247
rect 33793 20213 33827 20247
rect 34253 20213 34287 20247
rect 7757 20009 7791 20043
rect 19441 20009 19475 20043
rect 20545 20009 20579 20043
rect 23673 20009 23707 20043
rect 23765 20009 23799 20043
rect 28273 20009 28307 20043
rect 29561 20009 29595 20043
rect 31493 20009 31527 20043
rect 32781 20009 32815 20043
rect 34897 20009 34931 20043
rect 15761 19941 15795 19975
rect 26893 19941 26927 19975
rect 35449 19941 35483 19975
rect 7941 19873 7975 19907
rect 8033 19873 8067 19907
rect 8401 19873 8435 19907
rect 9505 19873 9539 19907
rect 12357 19873 12391 19907
rect 12449 19873 12483 19907
rect 12633 19873 12667 19907
rect 16221 19873 16255 19907
rect 16497 19873 16531 19907
rect 17877 19873 17911 19907
rect 18153 19873 18187 19907
rect 21005 19873 21039 19907
rect 23857 19873 23891 19907
rect 24777 19873 24811 19907
rect 32873 19873 32907 19907
rect 35541 19873 35575 19907
rect 8309 19805 8343 19839
rect 9229 19805 9263 19839
rect 10793 19805 10827 19839
rect 10885 19805 10919 19839
rect 10977 19802 11011 19836
rect 11137 19805 11171 19839
rect 12541 19805 12575 19839
rect 13369 19805 13403 19839
rect 14381 19805 14415 19839
rect 19993 19805 20027 19839
rect 20361 19805 20395 19839
rect 21281 19805 21315 19839
rect 22477 19805 22511 19839
rect 22845 19805 22879 19839
rect 23581 19805 23615 19839
rect 24593 19805 24627 19839
rect 24685 19805 24719 19839
rect 24869 19805 24903 19839
rect 25053 19805 25087 19839
rect 26065 19805 26099 19839
rect 26249 19805 26283 19839
rect 27169 19805 27203 19839
rect 29561 19805 29595 19839
rect 29745 19805 29779 19839
rect 30573 19805 30607 19839
rect 30757 19805 30791 19839
rect 31493 19805 31527 19839
rect 31677 19805 31711 19839
rect 32597 19805 32631 19839
rect 35078 19805 35112 19839
rect 14626 19737 14660 19771
rect 19349 19737 19383 19771
rect 20177 19737 20211 19771
rect 20269 19737 20303 19771
rect 22661 19737 22695 19771
rect 22753 19737 22787 19771
rect 26893 19737 26927 19771
rect 28089 19737 28123 19771
rect 28305 19737 28339 19771
rect 8217 19669 8251 19703
rect 10517 19669 10551 19703
rect 12173 19669 12207 19703
rect 13461 19669 13495 19703
rect 22017 19669 22051 19703
rect 23029 19669 23063 19703
rect 24409 19669 24443 19703
rect 26433 19669 26467 19703
rect 27077 19669 27111 19703
rect 28457 19669 28491 19703
rect 30757 19669 30791 19703
rect 32413 19669 32447 19703
rect 35081 19669 35115 19703
rect 9137 19465 9171 19499
rect 10149 19465 10183 19499
rect 14295 19465 14329 19499
rect 15485 19465 15519 19499
rect 18337 19465 18371 19499
rect 19441 19465 19475 19499
rect 20453 19465 20487 19499
rect 23029 19465 23063 19499
rect 25605 19465 25639 19499
rect 33885 19465 33919 19499
rect 35265 19465 35299 19499
rect 11621 19397 11655 19431
rect 11805 19397 11839 19431
rect 12633 19397 12667 19431
rect 14197 19397 14231 19431
rect 19165 19397 19199 19431
rect 20177 19397 20211 19431
rect 25881 19397 25915 19431
rect 26111 19397 26145 19431
rect 29653 19397 29687 19431
rect 29745 19397 29779 19431
rect 30665 19397 30699 19431
rect 30849 19397 30883 19431
rect 7757 19329 7791 19363
rect 8024 19329 8058 19363
rect 10333 19329 10367 19363
rect 10517 19329 10551 19363
rect 13461 19329 13495 19363
rect 13645 19329 13679 19363
rect 13737 19329 13771 19363
rect 14381 19329 14415 19363
rect 14473 19329 14507 19363
rect 15393 19329 15427 19363
rect 16957 19329 16991 19363
rect 17224 19329 17258 19363
rect 18889 19329 18923 19363
rect 19073 19329 19107 19363
rect 19257 19329 19291 19363
rect 19901 19329 19935 19363
rect 20085 19329 20119 19363
rect 20269 19329 20303 19363
rect 21005 19329 21039 19363
rect 22293 19329 22327 19363
rect 24041 19329 24075 19363
rect 25789 19329 25823 19363
rect 25973 19329 26007 19363
rect 26249 19329 26283 19363
rect 27537 19329 27571 19363
rect 28549 19329 28583 19363
rect 29561 19329 29595 19363
rect 29863 19329 29897 19363
rect 32137 19329 32171 19363
rect 32321 19329 32355 19363
rect 33021 19329 33055 19363
rect 33149 19329 33183 19363
rect 33241 19329 33275 19363
rect 34069 19329 34103 19363
rect 34161 19329 34195 19363
rect 34437 19329 34471 19363
rect 34897 19329 34931 19363
rect 10609 19261 10643 19295
rect 12265 19261 12299 19295
rect 15669 19261 15703 19295
rect 22017 19261 22051 19295
rect 24317 19261 24351 19295
rect 27813 19261 27847 19295
rect 28641 19261 28675 19295
rect 28917 19261 28951 19295
rect 30021 19261 30055 19295
rect 34989 19261 35023 19295
rect 12817 19193 12851 19227
rect 27629 19193 27663 19227
rect 34345 19193 34379 19227
rect 12633 19125 12667 19159
rect 13277 19125 13311 19159
rect 15025 19125 15059 19159
rect 21097 19125 21131 19159
rect 27721 19125 27755 19159
rect 29377 19125 29411 19159
rect 31033 19125 31067 19159
rect 32137 19125 32171 19159
rect 33425 19125 33459 19159
rect 35081 19125 35115 19159
rect 8125 18921 8159 18955
rect 9597 18921 9631 18955
rect 11253 18921 11287 18955
rect 13553 18921 13587 18955
rect 15761 18921 15795 18955
rect 21005 18921 21039 18955
rect 23673 18921 23707 18955
rect 23857 18921 23891 18955
rect 26157 18921 26191 18955
rect 28181 18921 28215 18955
rect 29561 18921 29595 18955
rect 30665 18921 30699 18955
rect 31769 18921 31803 18955
rect 24777 18853 24811 18887
rect 35265 18853 35299 18887
rect 10241 18785 10275 18819
rect 11621 18785 11655 18819
rect 23765 18785 23799 18819
rect 34989 18785 35023 18819
rect 8309 18717 8343 18751
rect 9505 18717 9539 18751
rect 9689 18717 9723 18751
rect 10333 18717 10367 18751
rect 11161 18717 11195 18751
rect 12173 18717 12207 18751
rect 14381 18717 14415 18751
rect 16405 18717 16439 18751
rect 16865 18717 16899 18751
rect 17877 18717 17911 18751
rect 18061 18717 18095 18751
rect 18245 18717 18279 18751
rect 19717 18717 19751 18751
rect 21925 18717 21959 18751
rect 22201 18717 22235 18751
rect 23581 18717 23615 18751
rect 24593 18717 24627 18751
rect 24685 18717 24719 18751
rect 24869 18717 24903 18751
rect 25053 18717 25087 18751
rect 25513 18717 25547 18751
rect 25881 18717 25915 18751
rect 25973 18717 26007 18751
rect 26617 18717 26651 18751
rect 26801 18717 26835 18751
rect 27077 18717 27111 18751
rect 28089 18717 28123 18751
rect 29745 18717 29779 18751
rect 29929 18717 29963 18751
rect 30205 18717 30239 18751
rect 30849 18717 30883 18751
rect 31125 18717 31159 18751
rect 31769 18717 31803 18751
rect 31861 18717 31895 18751
rect 32689 18717 32723 18751
rect 33057 18717 33091 18751
rect 33149 18717 33183 18751
rect 33333 18717 33367 18751
rect 33793 18717 33827 18751
rect 33977 18717 34011 18751
rect 34897 18717 34931 18751
rect 12440 18649 12474 18683
rect 14648 18649 14682 18683
rect 16221 18649 16255 18683
rect 16497 18649 16531 18683
rect 16589 18649 16623 18683
rect 16727 18649 16761 18683
rect 18153 18649 18187 18683
rect 23397 18649 23431 18683
rect 29837 18649 29871 18683
rect 30067 18649 30101 18683
rect 10701 18581 10735 18615
rect 18429 18581 18463 18615
rect 22937 18581 22971 18615
rect 24409 18581 24443 18615
rect 26985 18581 27019 18615
rect 28549 18581 28583 18615
rect 31033 18581 31067 18615
rect 32137 18581 32171 18615
rect 33885 18581 33919 18615
rect 12725 18377 12759 18411
rect 14013 18377 14047 18411
rect 16129 18377 16163 18411
rect 18061 18377 18095 18411
rect 21005 18377 21039 18411
rect 23765 18377 23799 18411
rect 25605 18377 25639 18411
rect 26249 18377 26283 18411
rect 29193 18377 29227 18411
rect 32505 18377 32539 18411
rect 33333 18377 33367 18411
rect 34989 18377 35023 18411
rect 9680 18309 9714 18343
rect 11989 18309 12023 18343
rect 12173 18309 12207 18343
rect 13921 18309 13955 18343
rect 15945 18309 15979 18343
rect 17049 18309 17083 18343
rect 17141 18309 17175 18343
rect 17969 18309 18003 18343
rect 26341 18309 26375 18343
rect 33149 18309 33183 18343
rect 9413 18241 9447 18275
rect 12909 18241 12943 18275
rect 13185 18241 13219 18275
rect 13369 18241 13403 18275
rect 15117 18241 15151 18275
rect 15301 18241 15335 18275
rect 15761 18241 15795 18275
rect 16865 18241 16899 18275
rect 17233 18241 17267 18275
rect 18705 18241 18739 18275
rect 18981 18241 19015 18275
rect 19993 18241 20027 18275
rect 20267 18241 20301 18275
rect 21833 18241 21867 18275
rect 22017 18241 22051 18275
rect 23029 18241 23063 18275
rect 24409 18241 24443 18275
rect 25513 18241 25547 18275
rect 25697 18241 25731 18275
rect 26157 18241 26191 18275
rect 26433 18241 26467 18275
rect 27905 18241 27939 18275
rect 28733 18241 28767 18275
rect 30849 18241 30883 18275
rect 32137 18241 32171 18275
rect 32965 18241 32999 18275
rect 33977 18241 34011 18275
rect 34805 18241 34839 18275
rect 34989 18241 35023 18275
rect 15209 18173 15243 18207
rect 22753 18173 22787 18207
rect 27997 18173 28031 18207
rect 30757 18173 30791 18207
rect 32229 18173 32263 18207
rect 34069 18173 34103 18207
rect 34345 18173 34379 18207
rect 10793 18105 10827 18139
rect 17417 18105 17451 18139
rect 31217 18105 31251 18139
rect 21833 18037 21867 18071
rect 24225 18037 24259 18071
rect 28181 18037 28215 18071
rect 28917 18037 28951 18071
rect 32137 18037 32171 18071
rect 10609 17833 10643 17867
rect 11345 17833 11379 17867
rect 14289 17833 14323 17867
rect 24593 17833 24627 17867
rect 24777 17833 24811 17867
rect 27721 17833 27755 17867
rect 30665 17833 30699 17867
rect 31401 17833 31435 17867
rect 18613 17765 18647 17799
rect 20269 17765 20303 17799
rect 21005 17765 21039 17799
rect 23581 17765 23615 17799
rect 25881 17765 25915 17799
rect 32321 17765 32355 17799
rect 15393 17697 15427 17731
rect 15577 17697 15611 17731
rect 16221 17697 16255 17731
rect 16497 17697 16531 17731
rect 17509 17697 17543 17731
rect 27261 17697 27295 17731
rect 10609 17629 10643 17663
rect 10793 17629 10827 17663
rect 11253 17629 11287 17663
rect 11437 17629 11471 17663
rect 14473 17629 14507 17663
rect 17693 17629 17727 17663
rect 18429 17629 18463 17663
rect 19257 17629 19291 17663
rect 19533 17629 19567 17663
rect 20821 17629 20855 17663
rect 20913 17629 20947 17663
rect 21557 17629 21591 17663
rect 21833 17629 21867 17663
rect 23029 17629 23063 17663
rect 23305 17629 23339 17663
rect 23397 17629 23431 17663
rect 25881 17629 25915 17663
rect 26157 17629 26191 17663
rect 27353 17629 27387 17663
rect 30573 17629 30607 17663
rect 30849 17629 30883 17663
rect 31309 17629 31343 17663
rect 31493 17629 31527 17663
rect 32229 17629 32263 17663
rect 32413 17629 32447 17663
rect 15301 17561 15335 17595
rect 23213 17561 23247 17595
rect 24409 17561 24443 17595
rect 30757 17561 30791 17595
rect 14933 17493 14967 17527
rect 17877 17493 17911 17527
rect 22569 17493 22603 17527
rect 24619 17493 24653 17527
rect 26065 17493 26099 17527
rect 12357 17289 12391 17323
rect 15577 17289 15611 17323
rect 21189 17289 21223 17323
rect 25973 17289 26007 17323
rect 10425 17221 10459 17255
rect 13737 17221 13771 17255
rect 16865 17221 16899 17255
rect 16957 17221 16991 17255
rect 17693 17221 17727 17255
rect 17909 17221 17943 17255
rect 20269 17221 20303 17255
rect 20361 17221 20395 17255
rect 10241 17153 10275 17187
rect 12541 17153 12575 17187
rect 12633 17153 12667 17187
rect 12909 17153 12943 17187
rect 13553 17153 13587 17187
rect 14464 17153 14498 17187
rect 16681 17153 16715 17187
rect 17049 17153 17083 17187
rect 19073 17153 19107 17187
rect 19257 17153 19291 17187
rect 19349 17153 19383 17187
rect 19441 17153 19475 17187
rect 20085 17153 20119 17187
rect 20453 17153 20487 17187
rect 21097 17153 21131 17187
rect 22109 17153 22143 17187
rect 23489 17153 23523 17187
rect 23765 17153 23799 17187
rect 24961 17153 24995 17187
rect 25237 17153 25271 17187
rect 13369 17085 13403 17119
rect 14197 17085 14231 17119
rect 21833 17085 21867 17119
rect 18061 17017 18095 17051
rect 12817 16949 12851 16983
rect 17233 16949 17267 16983
rect 17877 16949 17911 16983
rect 19625 16949 19659 16983
rect 20637 16949 20671 16983
rect 22845 16949 22879 16983
rect 24501 16949 24535 16983
rect 12357 16745 12391 16779
rect 12817 16745 12851 16779
rect 14105 16677 14139 16711
rect 14749 16677 14783 16711
rect 16865 16677 16899 16711
rect 18061 16677 18095 16711
rect 20361 16677 20395 16711
rect 9873 16609 9907 16643
rect 15485 16609 15519 16643
rect 25145 16609 25179 16643
rect 12541 16541 12575 16575
rect 12633 16541 12667 16575
rect 12909 16541 12943 16575
rect 13553 16541 13587 16575
rect 14105 16541 14139 16575
rect 14289 16541 14323 16575
rect 14933 16541 14967 16575
rect 15752 16541 15786 16575
rect 17877 16541 17911 16575
rect 18705 16541 18739 16575
rect 19349 16541 19383 16575
rect 19625 16541 19659 16575
rect 21465 16541 21499 16575
rect 21741 16541 21775 16575
rect 23397 16541 23431 16575
rect 25421 16541 25455 16575
rect 10118 16473 10152 16507
rect 11253 16405 11287 16439
rect 13369 16405 13403 16439
rect 18521 16405 18555 16439
rect 22477 16405 22511 16439
rect 23213 16405 23247 16439
rect 26525 16405 26559 16439
rect 11989 16201 12023 16235
rect 13829 16201 13863 16235
rect 16497 16201 16531 16235
rect 18521 16201 18555 16235
rect 22845 16201 22879 16235
rect 24961 16201 24995 16235
rect 25513 16201 25547 16235
rect 12716 16133 12750 16167
rect 22753 16133 22787 16167
rect 23826 16133 23860 16167
rect 7941 16065 7975 16099
rect 8585 16065 8619 16099
rect 8852 16065 8886 16099
rect 12449 16065 12483 16099
rect 14473 16065 14507 16099
rect 14740 16065 14774 16099
rect 17325 16065 17359 16099
rect 17785 16065 17819 16099
rect 18705 16065 18739 16099
rect 19441 16065 19475 16099
rect 20269 16065 20303 16099
rect 23581 16065 23615 16099
rect 25421 16065 25455 16099
rect 25605 16065 25639 16099
rect 26065 16065 26099 16099
rect 26249 16065 26283 16099
rect 11529 15997 11563 16031
rect 16037 15997 16071 16031
rect 17969 15997 18003 16031
rect 19993 15997 20027 16031
rect 22937 15997 22971 16031
rect 11805 15929 11839 15963
rect 15853 15929 15887 15963
rect 16313 15929 16347 15963
rect 19257 15929 19291 15963
rect 7757 15861 7791 15895
rect 9965 15861 9999 15895
rect 17601 15861 17635 15895
rect 21005 15861 21039 15895
rect 22385 15861 22419 15895
rect 26065 15861 26099 15895
rect 8953 15657 8987 15691
rect 9597 15657 9631 15691
rect 12541 15657 12575 15691
rect 13369 15657 13403 15691
rect 23765 15657 23799 15691
rect 25053 15657 25087 15691
rect 25973 15657 26007 15691
rect 12357 15589 12391 15623
rect 7021 15521 7055 15555
rect 9965 15521 9999 15555
rect 10057 15521 10091 15555
rect 10609 15521 10643 15555
rect 12081 15521 12115 15555
rect 13001 15521 13035 15555
rect 17693 15521 17727 15555
rect 19257 15521 19291 15555
rect 20729 15521 20763 15555
rect 22661 15521 22695 15555
rect 22845 15521 22879 15555
rect 26157 15521 26191 15555
rect 7288 15453 7322 15487
rect 9137 15453 9171 15487
rect 9781 15453 9815 15487
rect 9873 15453 9907 15487
rect 10885 15453 10919 15487
rect 10977 15453 11011 15487
rect 11069 15453 11103 15487
rect 11253 15453 11287 15487
rect 13185 15453 13219 15487
rect 15577 15453 15611 15487
rect 17969 15453 18003 15487
rect 19533 15453 19567 15487
rect 21005 15453 21039 15487
rect 23397 15453 23431 15487
rect 23581 15453 23615 15487
rect 24961 15453 24995 15487
rect 25881 15453 25915 15487
rect 15844 15385 15878 15419
rect 8401 15317 8435 15351
rect 16957 15317 16991 15351
rect 18705 15317 18739 15351
rect 20269 15317 20303 15351
rect 21741 15317 21775 15351
rect 22201 15317 22235 15351
rect 22569 15317 22603 15351
rect 25421 15317 25455 15351
rect 26157 15317 26191 15351
rect 8309 15113 8343 15147
rect 9137 15113 9171 15147
rect 12541 15113 12575 15147
rect 16681 15113 16715 15147
rect 21925 15113 21959 15147
rect 23949 15113 23983 15147
rect 7481 15045 7515 15079
rect 13430 15045 13464 15079
rect 21005 15045 21039 15079
rect 22814 15045 22848 15079
rect 6653 14977 6687 15011
rect 7297 14977 7331 15011
rect 8125 14977 8159 15011
rect 8953 14977 8987 15011
rect 9597 14977 9631 15011
rect 9864 14977 9898 15011
rect 11621 14977 11655 15011
rect 11713 14977 11747 15011
rect 12725 14977 12759 15011
rect 16865 14977 16899 15011
rect 18153 14977 18187 15011
rect 18429 14977 18463 15011
rect 20269 14977 20303 15011
rect 22109 14977 22143 15011
rect 24685 14977 24719 15011
rect 25697 14977 25731 15011
rect 7113 14909 7147 14943
rect 7941 14909 7975 14943
rect 8769 14909 8803 14943
rect 13185 14909 13219 14943
rect 20085 14909 20119 14943
rect 22569 14909 22603 14943
rect 24961 14909 24995 14943
rect 25421 14909 25455 14943
rect 24869 14841 24903 14875
rect 6469 14773 6503 14807
rect 10977 14773 11011 14807
rect 11897 14773 11931 14807
rect 14565 14773 14599 14807
rect 19165 14773 19199 14807
rect 20453 14773 20487 14807
rect 21097 14773 21131 14807
rect 24501 14773 24535 14807
rect 9689 14569 9723 14603
rect 9873 14569 9907 14603
rect 10609 14569 10643 14603
rect 10793 14569 10827 14603
rect 13093 14569 13127 14603
rect 16405 14569 16439 14603
rect 18705 14569 18739 14603
rect 23121 14569 23155 14603
rect 6837 14433 6871 14467
rect 10425 14433 10459 14467
rect 14197 14433 14231 14467
rect 24869 14433 24903 14467
rect 25053 14433 25087 14467
rect 25973 14433 26007 14467
rect 7093 14365 7127 14399
rect 10609 14365 10643 14399
rect 11713 14365 11747 14399
rect 11969 14365 12003 14399
rect 14381 14365 14415 14399
rect 15014 14365 15048 14399
rect 17325 14365 17359 14399
rect 19441 14365 19475 14399
rect 20085 14365 20119 14399
rect 21925 14365 21959 14399
rect 22109 14365 22143 14399
rect 22753 14365 22787 14399
rect 22937 14365 22971 14399
rect 23581 14365 23615 14399
rect 24777 14365 24811 14399
rect 26240 14365 26274 14399
rect 9505 14297 9539 14331
rect 10333 14297 10367 14331
rect 15292 14297 15326 14331
rect 17592 14297 17626 14331
rect 20330 14297 20364 14331
rect 8217 14229 8251 14263
rect 9715 14229 9749 14263
rect 14565 14229 14599 14263
rect 19257 14229 19291 14263
rect 21465 14229 21499 14263
rect 22293 14229 22327 14263
rect 23765 14229 23799 14263
rect 24409 14229 24443 14263
rect 27353 14229 27387 14263
rect 9965 14025 9999 14059
rect 11529 14025 11563 14059
rect 13645 14025 13679 14059
rect 18981 14025 19015 14059
rect 19717 14025 19751 14059
rect 20361 14025 20395 14059
rect 20729 14025 20763 14059
rect 22017 14025 22051 14059
rect 22477 14025 22511 14059
rect 25421 14025 25455 14059
rect 9781 13957 9815 13991
rect 12449 13957 12483 13991
rect 18889 13957 18923 13991
rect 20821 13957 20855 13991
rect 25237 13957 25271 13991
rect 25881 13957 25915 13991
rect 26081 13957 26115 13991
rect 28181 13957 28215 13991
rect 7941 13889 7975 13923
rect 8769 13889 8803 13923
rect 9413 13889 9447 13923
rect 9597 13889 9631 13923
rect 9689 13889 9723 13923
rect 10609 13889 10643 13923
rect 11713 13889 11747 13923
rect 12265 13889 12299 13923
rect 13461 13889 13495 13923
rect 15117 13889 15151 13923
rect 15209 13889 15243 13923
rect 15301 13889 15335 13923
rect 15485 13889 15519 13923
rect 16129 13889 16163 13923
rect 17049 13889 17083 13923
rect 17325 13889 17359 13923
rect 19901 13889 19935 13923
rect 22385 13889 22419 13923
rect 24133 13889 24167 13923
rect 27445 13889 27479 13923
rect 28089 13889 28123 13923
rect 7757 13821 7791 13855
rect 8125 13821 8159 13855
rect 8585 13821 8619 13855
rect 8953 13821 8987 13855
rect 13277 13821 13311 13855
rect 19073 13821 19107 13855
rect 20913 13821 20947 13855
rect 22569 13821 22603 13855
rect 23765 13821 23799 13855
rect 24225 13821 24259 13855
rect 24869 13821 24903 13855
rect 10425 13753 10459 13787
rect 27629 13753 27663 13787
rect 14841 13685 14875 13719
rect 15945 13685 15979 13719
rect 18521 13685 18555 13719
rect 24409 13685 24443 13719
rect 25237 13685 25271 13719
rect 26065 13685 26099 13719
rect 26249 13685 26283 13719
rect 8401 13481 8435 13515
rect 9689 13481 9723 13515
rect 10149 13481 10183 13515
rect 14473 13413 14507 13447
rect 18245 13413 18279 13447
rect 26525 13413 26559 13447
rect 7021 13345 7055 13379
rect 9781 13345 9815 13379
rect 13553 13345 13587 13379
rect 14841 13345 14875 13379
rect 15485 13345 15519 13379
rect 17877 13345 17911 13379
rect 19257 13345 19291 13379
rect 25053 13345 25087 13379
rect 25789 13345 25823 13379
rect 27261 13345 27295 13379
rect 9137 13277 9171 13311
rect 9965 13277 9999 13311
rect 11621 13277 11655 13311
rect 12725 13277 12759 13311
rect 13277 13277 13311 13311
rect 13369 13277 13403 13311
rect 14657 13277 14691 13311
rect 14749 13277 14783 13311
rect 14926 13277 14960 13311
rect 15752 13277 15786 13311
rect 18061 13277 18095 13311
rect 19441 13277 19475 13311
rect 21005 13277 21039 13311
rect 21465 13277 21499 13311
rect 23673 13277 23707 13311
rect 24869 13277 24903 13311
rect 25881 13277 25915 13311
rect 27537 13277 27571 13311
rect 7288 13209 7322 13243
rect 9689 13209 9723 13243
rect 11805 13209 11839 13243
rect 19625 13209 19659 13243
rect 21710 13209 21744 13243
rect 23857 13209 23891 13243
rect 25973 13209 26007 13243
rect 26341 13209 26375 13243
rect 8953 13141 8987 13175
rect 12541 13141 12575 13175
rect 16865 13141 16899 13175
rect 20821 13141 20855 13175
rect 22845 13141 22879 13175
rect 24409 13141 24443 13175
rect 24777 13141 24811 13175
rect 15669 12937 15703 12971
rect 16681 12937 16715 12971
rect 20085 12937 20119 12971
rect 22293 12937 22327 12971
rect 25789 12937 25823 12971
rect 13614 12869 13648 12903
rect 17570 12869 17604 12903
rect 27721 12869 27755 12903
rect 8033 12801 8067 12835
rect 8300 12801 8334 12835
rect 9965 12801 9999 12835
rect 10057 12801 10091 12835
rect 10977 12801 11011 12835
rect 11796 12801 11830 12835
rect 15209 12801 15243 12835
rect 15485 12801 15519 12835
rect 16865 12801 16899 12835
rect 19993 12801 20027 12835
rect 22201 12801 22235 12835
rect 23673 12801 23707 12835
rect 24133 12801 24167 12835
rect 24961 12801 24995 12835
rect 25053 12801 25087 12835
rect 25973 12801 26007 12835
rect 26065 12801 26099 12835
rect 26157 12801 26191 12835
rect 26341 12801 26375 12835
rect 26433 12801 26467 12835
rect 26985 12801 27019 12835
rect 27169 12801 27203 12835
rect 27537 12801 27571 12835
rect 28181 12801 28215 12835
rect 28365 12801 28399 12835
rect 37841 12801 37875 12835
rect 11529 12733 11563 12767
rect 13369 12733 13403 12767
rect 15393 12733 15427 12767
rect 17325 12733 17359 12767
rect 20177 12733 20211 12767
rect 22385 12733 22419 12767
rect 24869 12733 24903 12767
rect 25145 12733 25179 12767
rect 27261 12733 27295 12767
rect 27353 12733 27387 12767
rect 9413 12665 9447 12699
rect 10793 12665 10827 12699
rect 23489 12665 23523 12699
rect 28457 12665 28491 12699
rect 10241 12597 10275 12631
rect 12909 12597 12943 12631
rect 14749 12597 14783 12631
rect 15485 12597 15519 12631
rect 18705 12597 18739 12631
rect 19625 12597 19659 12631
rect 21833 12597 21867 12631
rect 24685 12597 24719 12631
rect 38025 12597 38059 12631
rect 8953 12393 8987 12427
rect 10977 12393 11011 12427
rect 13093 12393 13127 12427
rect 15117 12393 15151 12427
rect 15301 12393 15335 12427
rect 17233 12393 17267 12427
rect 17969 12393 18003 12427
rect 20637 12393 20671 12427
rect 27445 12393 27479 12427
rect 12633 12325 12667 12359
rect 9597 12257 9631 12291
rect 11437 12257 11471 12291
rect 12265 12257 12299 12291
rect 14105 12257 14139 12291
rect 16037 12257 16071 12291
rect 18429 12257 18463 12291
rect 18613 12257 18647 12291
rect 22385 12257 22419 12291
rect 23397 12257 23431 12291
rect 23489 12257 23523 12291
rect 24685 12257 24719 12291
rect 9137 12189 9171 12223
rect 11621 12189 11655 12223
rect 12449 12189 12483 12223
rect 13277 12189 13311 12223
rect 14289 12189 14323 12223
rect 15761 12189 15795 12223
rect 18337 12189 18371 12223
rect 19257 12189 19291 12223
rect 21281 12189 21315 12223
rect 22109 12189 22143 12223
rect 23305 12189 23339 12223
rect 24409 12189 24443 12223
rect 26249 12189 26283 12223
rect 26341 12189 26375 12223
rect 26525 12189 26559 12223
rect 26617 12189 26651 12223
rect 27077 12189 27111 12223
rect 27261 12189 27295 12223
rect 9842 12121 9876 12155
rect 11805 12121 11839 12155
rect 14933 12121 14967 12155
rect 17141 12121 17175 12155
rect 19524 12121 19558 12155
rect 26065 12121 26099 12155
rect 14473 12053 14507 12087
rect 15133 12053 15167 12087
rect 21097 12053 21131 12087
rect 21741 12053 21775 12087
rect 22201 12053 22235 12087
rect 22937 12053 22971 12087
rect 9505 11849 9539 11883
rect 14105 11849 14139 11883
rect 19533 11849 19567 11883
rect 27077 11849 27111 11883
rect 14994 11781 15028 11815
rect 8677 11713 8711 11747
rect 9689 11713 9723 11747
rect 10149 11713 10183 11747
rect 11529 11713 11563 11747
rect 13093 11713 13127 11747
rect 14289 11713 14323 11747
rect 14749 11713 14783 11747
rect 16957 11713 16991 11747
rect 18061 11713 18095 11747
rect 19349 11713 19383 11747
rect 20177 11713 20211 11747
rect 20361 11713 20395 11747
rect 21005 11713 21039 11747
rect 22937 11713 22971 11747
rect 23673 11713 23707 11747
rect 24961 11713 24995 11747
rect 25881 11713 25915 11747
rect 26985 11713 27019 11747
rect 27629 11713 27663 11747
rect 10425 11645 10459 11679
rect 12817 11645 12851 11679
rect 16681 11645 16715 11679
rect 19165 11645 19199 11679
rect 19993 11645 20027 11679
rect 22753 11645 22787 11679
rect 23949 11645 23983 11679
rect 25421 11645 25455 11679
rect 25973 11645 26007 11679
rect 27721 11645 27755 11679
rect 18245 11577 18279 11611
rect 8493 11509 8527 11543
rect 11713 11509 11747 11543
rect 16129 11509 16163 11543
rect 20821 11509 20855 11543
rect 23121 11509 23155 11543
rect 25053 11509 25087 11543
rect 25881 11509 25915 11543
rect 26249 11509 26283 11543
rect 12173 11305 12207 11339
rect 14749 11305 14783 11339
rect 24961 11305 24995 11339
rect 16313 11237 16347 11271
rect 18153 11237 18187 11271
rect 19257 11237 19291 11271
rect 22109 11237 22143 11271
rect 23857 11237 23891 11271
rect 26801 11237 26835 11271
rect 15485 11169 15519 11203
rect 15945 11169 15979 11203
rect 20729 11169 20763 11203
rect 1409 11101 1443 11135
rect 7021 11101 7055 11135
rect 8953 11101 8987 11135
rect 9209 11101 9243 11135
rect 10793 11101 10827 11135
rect 13277 11101 13311 11135
rect 13369 11101 13403 11135
rect 13553 11101 13587 11135
rect 14381 11101 14415 11135
rect 15301 11101 15335 11135
rect 16129 11101 16163 11135
rect 16773 11101 16807 11135
rect 19441 11101 19475 11135
rect 20985 11101 21019 11135
rect 23489 11101 23523 11135
rect 23673 11101 23707 11135
rect 24409 11101 24443 11135
rect 24782 11101 24816 11135
rect 25789 11101 25823 11135
rect 26341 11101 26375 11135
rect 26433 11101 26467 11135
rect 26709 11101 26743 11135
rect 26801 11101 26835 11135
rect 7288 11033 7322 11067
rect 11060 11033 11094 11067
rect 14197 11033 14231 11067
rect 17018 11033 17052 11067
rect 24593 11033 24627 11067
rect 24685 11033 24719 11067
rect 1593 10965 1627 10999
rect 8401 10965 8435 10999
rect 10333 10965 10367 10999
rect 14473 10965 14507 10999
rect 14565 10965 14599 10999
rect 7573 10761 7607 10795
rect 9689 10761 9723 10795
rect 10425 10761 10459 10795
rect 15393 10761 15427 10795
rect 15945 10761 15979 10795
rect 16865 10761 16899 10795
rect 19809 10761 19843 10795
rect 20729 10761 20763 10795
rect 8585 10693 8619 10727
rect 9229 10693 9263 10727
rect 14933 10693 14967 10727
rect 18061 10693 18095 10727
rect 18153 10693 18187 10727
rect 19441 10693 19475 10727
rect 19657 10693 19691 10727
rect 20269 10693 20303 10727
rect 24317 10693 24351 10727
rect 7757 10625 7791 10659
rect 8217 10625 8251 10659
rect 8401 10625 8435 10659
rect 9505 10625 9539 10659
rect 10793 10625 10827 10659
rect 11805 10625 11839 10659
rect 11897 10625 11931 10659
rect 11989 10625 12023 10659
rect 12173 10625 12207 10659
rect 13093 10625 13127 10659
rect 13360 10625 13394 10659
rect 15209 10625 15243 10659
rect 15853 10625 15887 10659
rect 17049 10625 17083 10659
rect 17785 10625 17819 10659
rect 17986 10615 18020 10649
rect 18271 10625 18305 10659
rect 20545 10625 20579 10659
rect 21833 10625 21867 10659
rect 22017 10625 22051 10659
rect 22845 10625 22879 10659
rect 26065 10625 26099 10659
rect 26341 10625 26375 10659
rect 9321 10557 9355 10591
rect 10609 10557 10643 10591
rect 10701 10557 10735 10591
rect 10885 10557 10919 10591
rect 11529 10557 11563 10591
rect 15025 10557 15059 10591
rect 17325 10557 17359 10591
rect 18429 10557 18463 10591
rect 20453 10557 20487 10591
rect 22661 10557 22695 10591
rect 24777 10557 24811 10591
rect 26249 10557 26283 10591
rect 24593 10489 24627 10523
rect 26161 10489 26195 10523
rect 9229 10421 9263 10455
rect 14473 10421 14507 10455
rect 14933 10421 14967 10455
rect 17233 10421 17267 10455
rect 19625 10421 19659 10455
rect 20269 10421 20303 10455
rect 22201 10421 22235 10455
rect 23029 10421 23063 10455
rect 25881 10421 25915 10455
rect 8401 10217 8435 10251
rect 10333 10217 10367 10251
rect 10517 10217 10551 10251
rect 14933 10217 14967 10251
rect 17049 10217 17083 10251
rect 17785 10217 17819 10251
rect 17969 10217 18003 10251
rect 20637 10217 20671 10251
rect 23029 10217 23063 10251
rect 24593 10217 24627 10251
rect 25421 10217 25455 10251
rect 24501 10149 24535 10183
rect 8033 10081 8067 10115
rect 15669 10081 15703 10115
rect 17693 10081 17727 10115
rect 21649 10081 21683 10115
rect 24685 10081 24719 10115
rect 8217 10013 8251 10047
rect 9321 10013 9355 10047
rect 9505 10013 9539 10047
rect 10977 10013 11011 10047
rect 12909 10013 12943 10047
rect 13001 10013 13035 10047
rect 14197 10013 14231 10047
rect 14289 10013 14323 10047
rect 15117 10013 15151 10047
rect 17509 10013 17543 10047
rect 17785 10013 17819 10047
rect 18613 10013 18647 10047
rect 19257 10013 19291 10047
rect 19513 10013 19547 10047
rect 24409 10013 24443 10047
rect 25329 10013 25363 10047
rect 25513 10013 25547 10047
rect 9137 9945 9171 9979
rect 10149 9945 10183 9979
rect 11222 9945 11256 9979
rect 13185 9945 13219 9979
rect 14473 9945 14507 9979
rect 15936 9945 15970 9979
rect 21916 9945 21950 9979
rect 9413 9877 9447 9911
rect 9689 9877 9723 9911
rect 10349 9877 10383 9911
rect 12357 9877 12391 9911
rect 18429 9877 18463 9911
rect 8585 9673 8619 9707
rect 10793 9673 10827 9707
rect 11989 9673 12023 9707
rect 15945 9673 15979 9707
rect 11529 9605 11563 9639
rect 17049 9605 17083 9639
rect 17960 9605 17994 9639
rect 7205 9537 7239 9571
rect 7472 9537 7506 9571
rect 9229 9537 9263 9571
rect 10977 9537 11011 9571
rect 11805 9537 11839 9571
rect 13369 9537 13403 9571
rect 13636 9537 13670 9571
rect 15393 9537 15427 9571
rect 16129 9537 16163 9571
rect 16865 9537 16899 9571
rect 17693 9537 17727 9571
rect 19901 9537 19935 9571
rect 20168 9537 20202 9571
rect 22201 9537 22235 9571
rect 22468 9537 22502 9571
rect 11621 9469 11655 9503
rect 16681 9469 16715 9503
rect 9045 9401 9079 9435
rect 15209 9401 15243 9435
rect 19073 9401 19107 9435
rect 11529 9333 11563 9367
rect 14749 9333 14783 9367
rect 21281 9333 21315 9367
rect 23581 9333 23615 9367
rect 8401 9129 8435 9163
rect 15485 9129 15519 9163
rect 18613 9129 18647 9163
rect 19625 9129 19659 9163
rect 21005 9129 21039 9163
rect 22109 9129 22143 9163
rect 22753 9129 22787 9163
rect 18061 9061 18095 9095
rect 8033 8993 8067 9027
rect 9505 8993 9539 9027
rect 12173 8993 12207 9027
rect 20177 8993 20211 9027
rect 8217 8925 8251 8959
rect 9689 8925 9723 8959
rect 10333 8925 10367 8959
rect 12357 8925 12391 8959
rect 13553 8925 13587 8959
rect 14105 8925 14139 8959
rect 16037 8925 16071 8959
rect 16129 8925 16163 8959
rect 16313 8925 16347 8959
rect 16957 8925 16991 8959
rect 18337 8925 18371 8959
rect 19257 8925 19291 8959
rect 19441 8925 19475 8959
rect 20361 8925 20395 8959
rect 20545 8925 20579 8959
rect 21189 8925 21223 8959
rect 22293 8925 22327 8959
rect 22937 8925 22971 8959
rect 10600 8857 10634 8891
rect 14350 8857 14384 8891
rect 18429 8857 18463 8891
rect 9873 8789 9907 8823
rect 11713 8789 11747 8823
rect 12541 8789 12575 8823
rect 13369 8789 13403 8823
rect 16773 8789 16807 8823
rect 18245 8789 18279 8823
rect 9597 8585 9631 8619
rect 10057 8585 10091 8619
rect 10701 8585 10735 8619
rect 13093 8585 13127 8619
rect 14197 8585 14231 8619
rect 16129 8585 16163 8619
rect 8484 8517 8518 8551
rect 15016 8517 15050 8551
rect 8217 8449 8251 8483
rect 10241 8449 10275 8483
rect 10885 8449 10919 8483
rect 11713 8449 11747 8483
rect 11980 8449 12014 8483
rect 13921 8449 13955 8483
rect 14013 8449 14047 8483
rect 17325 8449 17359 8483
rect 14749 8381 14783 8415
rect 17141 8245 17175 8279
rect 10885 8041 10919 8075
rect 11713 8041 11747 8075
rect 12173 8041 12207 8075
rect 18613 8041 18647 8075
rect 11345 7905 11379 7939
rect 17233 7905 17267 7939
rect 9505 7837 9539 7871
rect 11529 7837 11563 7871
rect 12357 7837 12391 7871
rect 17489 7837 17523 7871
rect 9772 7769 9806 7803
rect 9781 7497 9815 7531
rect 17601 7497 17635 7531
rect 9965 7361 9999 7395
rect 17233 7361 17267 7395
rect 17417 7361 17451 7395
rect 9045 6817 9079 6851
rect 9413 6817 9447 6851
rect 9229 6749 9263 6783
rect 1409 2601 1443 2635
rect 10425 2601 10459 2635
rect 31033 2465 31067 2499
rect 1593 2397 1627 2431
rect 10609 2397 10643 2431
rect 20729 2397 20763 2431
rect 30757 2397 30791 2431
rect 37841 2397 37875 2431
rect 20913 2261 20947 2295
rect 38025 2261 38059 2295
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 25222 37448 25228 37460
rect 25183 37420 25228 37448
rect 25222 37408 25228 37420
rect 25280 37408 25286 37460
rect 23845 37383 23903 37389
rect 23845 37349 23857 37383
rect 23891 37380 23903 37383
rect 24486 37380 24492 37392
rect 23891 37352 24492 37380
rect 23891 37349 23903 37352
rect 23845 37343 23903 37349
rect 24486 37340 24492 37352
rect 24544 37340 24550 37392
rect 25317 37383 25375 37389
rect 25317 37349 25329 37383
rect 25363 37380 25375 37383
rect 25498 37380 25504 37392
rect 25363 37352 25504 37380
rect 25363 37349 25375 37352
rect 25317 37343 25375 37349
rect 25498 37340 25504 37352
rect 25556 37340 25562 37392
rect 25866 37380 25872 37392
rect 25827 37352 25872 37380
rect 25866 37340 25872 37352
rect 25924 37340 25930 37392
rect 25225 37315 25283 37321
rect 25225 37281 25237 37315
rect 25271 37312 25283 37315
rect 27341 37315 27399 37321
rect 25271 37284 26372 37312
rect 25271 37281 25283 37284
rect 25225 37275 25283 37281
rect 3786 37244 3792 37256
rect 3747 37216 3792 37244
rect 3786 37204 3792 37216
rect 3844 37204 3850 37256
rect 14093 37247 14151 37253
rect 14093 37213 14105 37247
rect 14139 37244 14151 37247
rect 14918 37244 14924 37256
rect 14139 37216 14924 37244
rect 14139 37213 14151 37216
rect 14093 37207 14151 37213
rect 14918 37204 14924 37216
rect 14976 37204 14982 37256
rect 23661 37247 23719 37253
rect 23661 37213 23673 37247
rect 23707 37244 23719 37247
rect 23842 37244 23848 37256
rect 23707 37216 23848 37244
rect 23707 37213 23719 37216
rect 23661 37207 23719 37213
rect 23842 37204 23848 37216
rect 23900 37204 23906 37256
rect 25406 37244 25412 37256
rect 25367 37216 25412 37244
rect 25406 37204 25412 37216
rect 25464 37244 25470 37256
rect 26344 37253 26372 37284
rect 27341 37281 27353 37315
rect 27387 37312 27399 37315
rect 27614 37312 27620 37324
rect 27387 37284 27620 37312
rect 27387 37281 27399 37284
rect 27341 37275 27399 37281
rect 27614 37272 27620 37284
rect 27672 37312 27678 37324
rect 28537 37315 28595 37321
rect 28537 37312 28549 37315
rect 27672 37284 28549 37312
rect 27672 37272 27678 37284
rect 28537 37281 28549 37284
rect 28583 37281 28595 37315
rect 28537 37275 28595 37281
rect 26145 37247 26203 37253
rect 26145 37244 26157 37247
rect 25464 37216 26157 37244
rect 25464 37204 25470 37216
rect 26145 37213 26157 37216
rect 26191 37213 26203 37247
rect 26145 37207 26203 37213
rect 26329 37247 26387 37253
rect 26329 37213 26341 37247
rect 26375 37244 26387 37247
rect 26418 37244 26424 37256
rect 26375 37216 26424 37244
rect 26375 37213 26387 37216
rect 26329 37207 26387 37213
rect 26418 37204 26424 37216
rect 26476 37204 26482 37256
rect 28626 37244 28632 37256
rect 26896 37216 28396 37244
rect 28539 37216 28632 37244
rect 25041 37179 25099 37185
rect 25041 37145 25053 37179
rect 25087 37176 25099 37179
rect 26896 37176 26924 37216
rect 25087 37148 26924 37176
rect 25087 37145 25099 37148
rect 25041 37139 25099 37145
rect 26970 37136 26976 37188
rect 27028 37176 27034 37188
rect 27157 37179 27215 37185
rect 27028 37148 27073 37176
rect 27028 37136 27034 37148
rect 27157 37145 27169 37179
rect 27203 37145 27215 37179
rect 28258 37176 28264 37188
rect 28219 37148 28264 37176
rect 27157 37139 27215 37145
rect 3234 37068 3240 37120
rect 3292 37108 3298 37120
rect 3973 37111 4031 37117
rect 3973 37108 3985 37111
rect 3292 37080 3985 37108
rect 3292 37068 3298 37080
rect 3973 37077 3985 37080
rect 4019 37077 4031 37111
rect 3973 37071 4031 37077
rect 13538 37068 13544 37120
rect 13596 37108 13602 37120
rect 14277 37111 14335 37117
rect 14277 37108 14289 37111
rect 13596 37080 14289 37108
rect 13596 37068 13602 37080
rect 14277 37077 14289 37080
rect 14323 37077 14335 37111
rect 14277 37071 14335 37077
rect 26053 37111 26111 37117
rect 26053 37077 26065 37111
rect 26099 37108 26111 37111
rect 26326 37108 26332 37120
rect 26099 37080 26332 37108
rect 26099 37077 26111 37080
rect 26053 37071 26111 37077
rect 26326 37068 26332 37080
rect 26384 37068 26390 37120
rect 26418 37068 26424 37120
rect 26476 37108 26482 37120
rect 27172 37108 27200 37139
rect 28258 37136 28264 37148
rect 28316 37136 28322 37188
rect 28368 37176 28396 37216
rect 28626 37204 28632 37216
rect 28684 37244 28690 37256
rect 30282 37244 30288 37256
rect 28684 37216 30288 37244
rect 28684 37204 28690 37216
rect 30282 37204 30288 37216
rect 30340 37204 30346 37256
rect 30469 37247 30527 37253
rect 30469 37213 30481 37247
rect 30515 37213 30527 37247
rect 30469 37207 30527 37213
rect 34701 37247 34759 37253
rect 34701 37213 34713 37247
rect 34747 37244 34759 37247
rect 35802 37244 35808 37256
rect 34747 37216 35808 37244
rect 34747 37213 34759 37216
rect 34701 37207 34759 37213
rect 28721 37179 28779 37185
rect 28721 37176 28733 37179
rect 28368 37148 28733 37176
rect 28721 37145 28733 37148
rect 28767 37145 28779 37179
rect 28721 37139 28779 37145
rect 29730 37136 29736 37188
rect 29788 37176 29794 37188
rect 30484 37176 30512 37207
rect 35802 37204 35808 37216
rect 35860 37204 35866 37256
rect 29788 37148 30512 37176
rect 29788 37136 29794 37148
rect 26476 37080 27200 37108
rect 28353 37111 28411 37117
rect 26476 37068 26482 37080
rect 28353 37077 28365 37111
rect 28399 37108 28411 37111
rect 28810 37108 28816 37120
rect 28399 37080 28816 37108
rect 28399 37077 28411 37080
rect 28353 37071 28411 37077
rect 28810 37068 28816 37080
rect 28868 37068 28874 37120
rect 30377 37111 30435 37117
rect 30377 37077 30389 37111
rect 30423 37108 30435 37111
rect 30466 37108 30472 37120
rect 30423 37080 30472 37108
rect 30423 37077 30435 37080
rect 30377 37071 30435 37077
rect 30466 37068 30472 37080
rect 30524 37068 30530 37120
rect 34514 37068 34520 37120
rect 34572 37108 34578 37120
rect 34885 37111 34943 37117
rect 34885 37108 34897 37111
rect 34572 37080 34897 37108
rect 34572 37068 34578 37080
rect 34885 37077 34897 37080
rect 34931 37077 34943 37111
rect 34885 37071 34943 37077
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 25222 36864 25228 36916
rect 25280 36904 25286 36916
rect 25409 36907 25467 36913
rect 25409 36904 25421 36907
rect 25280 36876 25421 36904
rect 25280 36864 25286 36876
rect 25409 36873 25421 36876
rect 25455 36873 25467 36907
rect 28810 36904 28816 36916
rect 28771 36876 28816 36904
rect 25409 36867 25467 36873
rect 28810 36864 28816 36876
rect 28868 36904 28874 36916
rect 29638 36904 29644 36916
rect 28868 36876 29644 36904
rect 28868 36864 28874 36876
rect 29638 36864 29644 36876
rect 29696 36904 29702 36916
rect 29733 36907 29791 36913
rect 29733 36904 29745 36907
rect 29696 36876 29745 36904
rect 29696 36864 29702 36876
rect 29733 36873 29745 36876
rect 29779 36873 29791 36907
rect 29733 36867 29791 36873
rect 24394 36836 24400 36848
rect 24355 36808 24400 36836
rect 24394 36796 24400 36808
rect 24452 36796 24458 36848
rect 25317 36839 25375 36845
rect 25317 36805 25329 36839
rect 25363 36836 25375 36839
rect 26237 36839 26295 36845
rect 26237 36836 26249 36839
rect 25363 36808 26249 36836
rect 25363 36805 25375 36808
rect 25317 36799 25375 36805
rect 26237 36805 26249 36808
rect 26283 36805 26295 36839
rect 26237 36799 26295 36805
rect 28258 36796 28264 36848
rect 28316 36836 28322 36848
rect 28316 36808 28948 36836
rect 28316 36796 28322 36808
rect 24213 36771 24271 36777
rect 24213 36737 24225 36771
rect 24259 36768 24271 36771
rect 24302 36768 24308 36780
rect 24259 36740 24308 36768
rect 24259 36737 24271 36740
rect 24213 36731 24271 36737
rect 24302 36728 24308 36740
rect 24360 36728 24366 36780
rect 24489 36771 24547 36777
rect 24489 36737 24501 36771
rect 24535 36768 24547 36771
rect 24762 36768 24768 36780
rect 24535 36740 24768 36768
rect 24535 36737 24547 36740
rect 24489 36731 24547 36737
rect 24762 36728 24768 36740
rect 24820 36768 24826 36780
rect 26145 36771 26203 36777
rect 26145 36768 26157 36771
rect 24820 36740 26157 36768
rect 24820 36728 24826 36740
rect 26145 36737 26157 36740
rect 26191 36737 26203 36771
rect 26145 36731 26203 36737
rect 26329 36771 26387 36777
rect 26329 36737 26341 36771
rect 26375 36737 26387 36771
rect 26329 36731 26387 36737
rect 27433 36771 27491 36777
rect 27433 36737 27445 36771
rect 27479 36768 27491 36771
rect 27614 36768 27620 36780
rect 27479 36740 27620 36768
rect 27479 36737 27491 36740
rect 27433 36731 27491 36737
rect 25593 36703 25651 36709
rect 25593 36669 25605 36703
rect 25639 36669 25651 36703
rect 25593 36663 25651 36669
rect 24213 36635 24271 36641
rect 24213 36601 24225 36635
rect 24259 36632 24271 36635
rect 25498 36632 25504 36644
rect 24259 36604 25504 36632
rect 24259 36601 24271 36604
rect 24213 36595 24271 36601
rect 25498 36592 25504 36604
rect 25556 36592 25562 36644
rect 24946 36564 24952 36576
rect 24907 36536 24952 36564
rect 24946 36524 24952 36536
rect 25004 36524 25010 36576
rect 25608 36564 25636 36663
rect 26234 36660 26240 36712
rect 26292 36700 26298 36712
rect 26344 36700 26372 36731
rect 27614 36728 27620 36740
rect 27672 36728 27678 36780
rect 28626 36768 28632 36780
rect 28587 36740 28632 36768
rect 28626 36728 28632 36740
rect 28684 36728 28690 36780
rect 28920 36777 28948 36808
rect 28905 36771 28963 36777
rect 28905 36737 28917 36771
rect 28951 36737 28963 36771
rect 28905 36731 28963 36737
rect 29641 36771 29699 36777
rect 29641 36737 29653 36771
rect 29687 36768 29699 36771
rect 29730 36768 29736 36780
rect 29687 36740 29736 36768
rect 29687 36737 29699 36740
rect 29641 36731 29699 36737
rect 26292 36672 26372 36700
rect 27525 36703 27583 36709
rect 26292 36660 26298 36672
rect 27525 36669 27537 36703
rect 27571 36700 27583 36703
rect 28445 36703 28503 36709
rect 28445 36700 28457 36703
rect 27571 36672 28457 36700
rect 27571 36669 27583 36672
rect 27525 36663 27583 36669
rect 28445 36669 28457 36672
rect 28491 36669 28503 36703
rect 28920 36700 28948 36731
rect 29730 36728 29736 36740
rect 29788 36728 29794 36780
rect 29822 36728 29828 36780
rect 29880 36768 29886 36780
rect 30466 36768 30472 36780
rect 29880 36740 29925 36768
rect 30427 36740 30472 36768
rect 29880 36728 29886 36740
rect 30466 36728 30472 36740
rect 30524 36728 30530 36780
rect 30190 36700 30196 36712
rect 28920 36672 30196 36700
rect 28445 36663 28503 36669
rect 30190 36660 30196 36672
rect 30248 36700 30254 36712
rect 30561 36703 30619 36709
rect 30248 36672 30512 36700
rect 30248 36660 30254 36672
rect 26326 36592 26332 36644
rect 26384 36632 26390 36644
rect 30374 36632 30380 36644
rect 26384 36604 30380 36632
rect 26384 36592 26390 36604
rect 30374 36592 30380 36604
rect 30432 36592 30438 36644
rect 30484 36632 30512 36672
rect 30561 36669 30573 36703
rect 30607 36700 30619 36703
rect 30926 36700 30932 36712
rect 30607 36672 30932 36700
rect 30607 36669 30619 36672
rect 30561 36663 30619 36669
rect 30926 36660 30932 36672
rect 30984 36660 30990 36712
rect 32490 36632 32496 36644
rect 30484 36604 32496 36632
rect 32490 36592 32496 36604
rect 32548 36592 32554 36644
rect 27522 36564 27528 36576
rect 25608 36536 27528 36564
rect 27522 36524 27528 36536
rect 27580 36524 27586 36576
rect 27706 36564 27712 36576
rect 27667 36536 27712 36564
rect 27706 36524 27712 36536
rect 27764 36524 27770 36576
rect 28902 36524 28908 36576
rect 28960 36564 28966 36576
rect 30745 36567 30803 36573
rect 30745 36564 30757 36567
rect 28960 36536 30757 36564
rect 28960 36524 28966 36536
rect 30745 36533 30757 36536
rect 30791 36533 30803 36567
rect 30745 36527 30803 36533
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 23753 36363 23811 36369
rect 23753 36329 23765 36363
rect 23799 36360 23811 36363
rect 24394 36360 24400 36372
rect 23799 36332 24400 36360
rect 23799 36329 23811 36332
rect 23753 36323 23811 36329
rect 24394 36320 24400 36332
rect 24452 36360 24458 36372
rect 24949 36363 25007 36369
rect 24949 36360 24961 36363
rect 24452 36332 24961 36360
rect 24452 36320 24458 36332
rect 24949 36329 24961 36332
rect 24995 36360 25007 36363
rect 26050 36360 26056 36372
rect 24995 36332 26056 36360
rect 24995 36329 25007 36332
rect 24949 36323 25007 36329
rect 26050 36320 26056 36332
rect 26108 36320 26114 36372
rect 26234 36360 26240 36372
rect 26195 36332 26240 36360
rect 26234 36320 26240 36332
rect 26292 36360 26298 36372
rect 26970 36360 26976 36372
rect 26292 36332 26976 36360
rect 26292 36320 26298 36332
rect 26970 36320 26976 36332
rect 27028 36320 27034 36372
rect 27522 36320 27528 36372
rect 27580 36360 27586 36372
rect 28810 36360 28816 36372
rect 27580 36332 28816 36360
rect 27580 36320 27586 36332
rect 28810 36320 28816 36332
rect 28868 36320 28874 36372
rect 29825 36363 29883 36369
rect 29825 36329 29837 36363
rect 29871 36360 29883 36363
rect 30653 36363 30711 36369
rect 29871 36332 30144 36360
rect 29871 36329 29883 36332
rect 29825 36323 29883 36329
rect 25133 36295 25191 36301
rect 25133 36261 25145 36295
rect 25179 36292 25191 36295
rect 25406 36292 25412 36304
rect 25179 36264 25412 36292
rect 25179 36261 25191 36264
rect 25133 36255 25191 36261
rect 25406 36252 25412 36264
rect 25464 36292 25470 36304
rect 28902 36292 28908 36304
rect 25464 36264 26280 36292
rect 25464 36252 25470 36264
rect 26252 36233 26280 36264
rect 28736 36264 28908 36292
rect 28736 36233 28764 36264
rect 28902 36252 28908 36264
rect 28960 36252 28966 36304
rect 30009 36295 30067 36301
rect 30009 36261 30021 36295
rect 30055 36261 30067 36295
rect 30116 36292 30144 36332
rect 30653 36329 30665 36363
rect 30699 36360 30711 36363
rect 30926 36360 30932 36372
rect 30699 36332 30788 36360
rect 30887 36332 30932 36360
rect 30699 36329 30711 36332
rect 30653 36323 30711 36329
rect 30282 36292 30288 36304
rect 30116 36264 30288 36292
rect 30009 36255 30067 36261
rect 26237 36227 26295 36233
rect 26237 36193 26249 36227
rect 26283 36193 26295 36227
rect 26237 36187 26295 36193
rect 28721 36227 28779 36233
rect 28721 36193 28733 36227
rect 28767 36193 28779 36227
rect 28721 36187 28779 36193
rect 28810 36184 28816 36236
rect 28868 36224 28874 36236
rect 30024 36224 30052 36255
rect 30282 36252 30288 36264
rect 30340 36292 30346 36304
rect 30760 36292 30788 36332
rect 30926 36320 30932 36332
rect 30984 36320 30990 36372
rect 31570 36360 31576 36372
rect 31531 36332 31576 36360
rect 31570 36320 31576 36332
rect 31628 36320 31634 36372
rect 30340 36264 30696 36292
rect 30760 36264 31708 36292
rect 30340 36252 30346 36264
rect 30668 36224 30696 36264
rect 31481 36227 31539 36233
rect 28868 36196 28913 36224
rect 30024 36196 30604 36224
rect 30668 36196 31432 36224
rect 28868 36184 28874 36196
rect 23661 36159 23719 36165
rect 23661 36125 23673 36159
rect 23707 36156 23719 36159
rect 25038 36156 25044 36168
rect 23707 36128 25044 36156
rect 23707 36125 23719 36128
rect 23661 36119 23719 36125
rect 25038 36116 25044 36128
rect 25096 36116 25102 36168
rect 25866 36116 25872 36168
rect 25924 36156 25930 36168
rect 26145 36159 26203 36165
rect 26145 36156 26157 36159
rect 25924 36128 26157 36156
rect 25924 36116 25930 36128
rect 26145 36125 26157 36128
rect 26191 36125 26203 36159
rect 26418 36156 26424 36168
rect 26379 36128 26424 36156
rect 26145 36119 26203 36125
rect 26418 36116 26424 36128
rect 26476 36116 26482 36168
rect 29638 36156 29644 36168
rect 29599 36128 29644 36156
rect 29638 36116 29644 36128
rect 29696 36116 29702 36168
rect 29733 36159 29791 36165
rect 29733 36125 29745 36159
rect 29779 36125 29791 36159
rect 29733 36119 29791 36125
rect 24302 36048 24308 36100
rect 24360 36088 24366 36100
rect 24765 36091 24823 36097
rect 24765 36088 24777 36091
rect 24360 36060 24777 36088
rect 24360 36048 24366 36060
rect 24765 36057 24777 36060
rect 24811 36057 24823 36091
rect 29748 36088 29776 36119
rect 30190 36116 30196 36168
rect 30248 36156 30254 36168
rect 30469 36159 30527 36165
rect 30469 36156 30481 36159
rect 30248 36128 30481 36156
rect 30248 36116 30254 36128
rect 30469 36125 30481 36128
rect 30515 36125 30527 36159
rect 30576 36156 30604 36196
rect 31202 36156 31208 36168
rect 30576 36128 31208 36156
rect 30469 36119 30527 36125
rect 31202 36116 31208 36128
rect 31260 36116 31266 36168
rect 31404 36165 31432 36196
rect 31481 36193 31493 36227
rect 31527 36193 31539 36227
rect 31481 36187 31539 36193
rect 31389 36159 31447 36165
rect 31389 36125 31401 36159
rect 31435 36125 31447 36159
rect 31389 36119 31447 36125
rect 31294 36088 31300 36100
rect 24765 36051 24823 36057
rect 26620 36060 31300 36088
rect 24854 35980 24860 36032
rect 24912 36020 24918 36032
rect 26620 36029 26648 36060
rect 31294 36048 31300 36060
rect 31352 36048 31358 36100
rect 31496 36088 31524 36187
rect 31680 36168 31708 36264
rect 32122 36184 32128 36236
rect 32180 36224 32186 36236
rect 32585 36227 32643 36233
rect 32585 36224 32597 36227
rect 32180 36196 32597 36224
rect 32180 36184 32186 36196
rect 32585 36193 32597 36196
rect 32631 36193 32643 36227
rect 32585 36187 32643 36193
rect 31662 36156 31668 36168
rect 31623 36128 31668 36156
rect 31662 36116 31668 36128
rect 31720 36116 31726 36168
rect 32214 36116 32220 36168
rect 32272 36156 32278 36168
rect 32309 36159 32367 36165
rect 32309 36156 32321 36159
rect 32272 36128 32321 36156
rect 32272 36116 32278 36128
rect 32309 36125 32321 36128
rect 32355 36125 32367 36159
rect 32309 36119 32367 36125
rect 32398 36116 32404 36168
rect 32456 36156 32462 36168
rect 32456 36128 32501 36156
rect 32456 36116 32462 36128
rect 31404 36060 31524 36088
rect 24965 36023 25023 36029
rect 24965 36020 24977 36023
rect 24912 35992 24977 36020
rect 24912 35980 24918 35992
rect 24965 35989 24977 35992
rect 25011 35989 25023 36023
rect 24965 35983 25023 35989
rect 26605 36023 26663 36029
rect 26605 35989 26617 36023
rect 26651 35989 26663 36023
rect 28258 36020 28264 36032
rect 28219 35992 28264 36020
rect 26605 35983 26663 35989
rect 28258 35980 28264 35992
rect 28316 35980 28322 36032
rect 28626 36020 28632 36032
rect 28587 35992 28632 36020
rect 28626 35980 28632 35992
rect 28684 35980 28690 36032
rect 30282 35980 30288 36032
rect 30340 36020 30346 36032
rect 31404 36020 31432 36060
rect 31846 36020 31852 36032
rect 30340 35992 31432 36020
rect 31807 35992 31852 36020
rect 30340 35980 30346 35992
rect 31846 35980 31852 35992
rect 31904 35980 31910 36032
rect 32585 36023 32643 36029
rect 32585 35989 32597 36023
rect 32631 36020 32643 36023
rect 32950 36020 32956 36032
rect 32631 35992 32956 36020
rect 32631 35989 32643 35992
rect 32585 35983 32643 35989
rect 32950 35980 32956 35992
rect 33008 35980 33014 36032
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 24762 35816 24768 35828
rect 24723 35788 24768 35816
rect 24762 35776 24768 35788
rect 24820 35776 24826 35828
rect 26142 35776 26148 35828
rect 26200 35816 26206 35828
rect 26329 35819 26387 35825
rect 26329 35816 26341 35819
rect 26200 35788 26341 35816
rect 26200 35776 26206 35788
rect 26329 35785 26341 35788
rect 26375 35785 26387 35819
rect 26329 35779 26387 35785
rect 27433 35819 27491 35825
rect 27433 35785 27445 35819
rect 27479 35816 27491 35819
rect 27706 35816 27712 35828
rect 27479 35788 27712 35816
rect 27479 35785 27491 35788
rect 27433 35779 27491 35785
rect 27706 35776 27712 35788
rect 27764 35776 27770 35828
rect 28534 35816 28540 35828
rect 28368 35788 28540 35816
rect 25961 35751 26019 35757
rect 25240 35720 25912 35748
rect 23569 35683 23627 35689
rect 23569 35649 23581 35683
rect 23615 35649 23627 35683
rect 23750 35680 23756 35692
rect 23711 35652 23756 35680
rect 23569 35643 23627 35649
rect 23584 35612 23612 35643
rect 23750 35640 23756 35652
rect 23808 35640 23814 35692
rect 24394 35640 24400 35692
rect 24452 35680 24458 35692
rect 25240 35689 25268 35720
rect 24949 35683 25007 35689
rect 24949 35680 24961 35683
rect 24452 35652 24961 35680
rect 24452 35640 24458 35652
rect 24949 35649 24961 35652
rect 24995 35649 25007 35683
rect 24949 35643 25007 35649
rect 25041 35683 25099 35689
rect 25041 35649 25053 35683
rect 25087 35649 25099 35683
rect 25041 35643 25099 35649
rect 25225 35683 25283 35689
rect 25225 35649 25237 35683
rect 25271 35649 25283 35683
rect 25225 35643 25283 35649
rect 24026 35612 24032 35624
rect 23584 35584 24032 35612
rect 24026 35572 24032 35584
rect 24084 35572 24090 35624
rect 25056 35612 25084 35643
rect 25314 35640 25320 35692
rect 25372 35680 25378 35692
rect 25372 35652 25417 35680
rect 25372 35640 25378 35652
rect 25406 35612 25412 35624
rect 25056 35584 25412 35612
rect 25406 35572 25412 35584
rect 25464 35572 25470 35624
rect 25884 35612 25912 35720
rect 25961 35717 25973 35751
rect 26007 35748 26019 35751
rect 27341 35751 27399 35757
rect 27341 35748 27353 35751
rect 26007 35720 27353 35748
rect 26007 35717 26019 35720
rect 25961 35711 26019 35717
rect 27341 35717 27353 35720
rect 27387 35717 27399 35751
rect 28368 35748 28396 35788
rect 28534 35776 28540 35788
rect 28592 35816 28598 35828
rect 29473 35819 29531 35825
rect 29473 35816 29485 35819
rect 28592 35788 29485 35816
rect 28592 35776 28598 35788
rect 29473 35785 29485 35788
rect 29519 35785 29531 35819
rect 29473 35779 29531 35785
rect 29641 35819 29699 35825
rect 29641 35785 29653 35819
rect 29687 35816 29699 35819
rect 29730 35816 29736 35828
rect 29687 35788 29736 35816
rect 29687 35785 29699 35788
rect 29641 35779 29699 35785
rect 29730 35776 29736 35788
rect 29788 35816 29794 35828
rect 30282 35816 30288 35828
rect 29788 35788 30288 35816
rect 29788 35776 29794 35788
rect 30282 35776 30288 35788
rect 30340 35776 30346 35828
rect 32490 35816 32496 35828
rect 32451 35788 32496 35816
rect 32490 35776 32496 35788
rect 32548 35776 32554 35828
rect 28718 35748 28724 35760
rect 27341 35711 27399 35717
rect 28276 35720 28396 35748
rect 28679 35720 28724 35748
rect 26145 35683 26203 35689
rect 26145 35649 26157 35683
rect 26191 35680 26203 35683
rect 26326 35680 26332 35692
rect 26191 35652 26332 35680
rect 26191 35649 26203 35652
rect 26145 35643 26203 35649
rect 26326 35640 26332 35652
rect 26384 35640 26390 35692
rect 26421 35683 26479 35689
rect 26421 35649 26433 35683
rect 26467 35680 26479 35683
rect 26786 35680 26792 35692
rect 26467 35652 26792 35680
rect 26467 35649 26479 35652
rect 26421 35643 26479 35649
rect 26786 35640 26792 35652
rect 26844 35640 26850 35692
rect 28276 35689 28304 35720
rect 28718 35708 28724 35720
rect 28776 35708 28782 35760
rect 29273 35751 29331 35757
rect 29273 35748 29285 35751
rect 28828 35720 29285 35748
rect 28261 35683 28319 35689
rect 28261 35649 28273 35683
rect 28307 35649 28319 35683
rect 28442 35680 28448 35692
rect 28403 35652 28448 35680
rect 28261 35643 28319 35649
rect 28442 35640 28448 35652
rect 28500 35640 28506 35692
rect 26510 35612 26516 35624
rect 25884 35584 26516 35612
rect 26510 35572 26516 35584
rect 26568 35572 26574 35624
rect 27522 35612 27528 35624
rect 27483 35584 27528 35612
rect 27522 35572 27528 35584
rect 27580 35572 27586 35624
rect 28350 35572 28356 35624
rect 28408 35612 28414 35624
rect 28828 35621 28856 35720
rect 29273 35717 29285 35720
rect 29319 35717 29331 35751
rect 32508 35748 32536 35776
rect 32508 35720 33180 35748
rect 29273 35711 29331 35717
rect 30374 35640 30380 35692
rect 30432 35680 30438 35692
rect 31113 35683 31171 35689
rect 31113 35680 31125 35683
rect 30432 35652 31125 35680
rect 30432 35640 30438 35652
rect 31113 35649 31125 35652
rect 31159 35649 31171 35683
rect 31294 35680 31300 35692
rect 31255 35652 31300 35680
rect 31113 35643 31171 35649
rect 31294 35640 31300 35652
rect 31352 35640 31358 35692
rect 31573 35683 31631 35689
rect 31573 35649 31585 35683
rect 31619 35680 31631 35683
rect 32122 35680 32128 35692
rect 31619 35652 31984 35680
rect 32083 35652 32128 35680
rect 31619 35649 31631 35652
rect 31573 35643 31631 35649
rect 28813 35615 28871 35621
rect 28813 35612 28825 35615
rect 28408 35584 28825 35612
rect 28408 35572 28414 35584
rect 28813 35581 28825 35584
rect 28859 35581 28871 35615
rect 28813 35575 28871 35581
rect 31205 35615 31263 35621
rect 31205 35581 31217 35615
rect 31251 35612 31263 35615
rect 31846 35612 31852 35624
rect 31251 35584 31852 35612
rect 31251 35581 31263 35584
rect 31205 35575 31263 35581
rect 31846 35572 31852 35584
rect 31904 35572 31910 35624
rect 31956 35612 31984 35652
rect 32122 35640 32128 35652
rect 32180 35640 32186 35692
rect 32950 35680 32956 35692
rect 32911 35652 32956 35680
rect 32950 35640 32956 35652
rect 33008 35640 33014 35692
rect 33152 35689 33180 35720
rect 33137 35683 33195 35689
rect 33137 35649 33149 35683
rect 33183 35649 33195 35683
rect 33137 35643 33195 35649
rect 32214 35612 32220 35624
rect 31956 35584 32220 35612
rect 32214 35572 32220 35584
rect 32272 35572 32278 35624
rect 23842 35504 23848 35556
rect 23900 35544 23906 35556
rect 28166 35544 28172 35556
rect 23900 35516 28172 35544
rect 23900 35504 23906 35516
rect 28166 35504 28172 35516
rect 28224 35504 28230 35556
rect 23658 35476 23664 35488
rect 23619 35448 23664 35476
rect 23658 35436 23664 35448
rect 23716 35436 23722 35488
rect 26973 35479 27031 35485
rect 26973 35445 26985 35479
rect 27019 35476 27031 35479
rect 27246 35476 27252 35488
rect 27019 35448 27252 35476
rect 27019 35445 27031 35448
rect 26973 35439 27031 35445
rect 27246 35436 27252 35448
rect 27304 35436 27310 35488
rect 28442 35436 28448 35488
rect 28500 35476 28506 35488
rect 29457 35479 29515 35485
rect 29457 35476 29469 35479
rect 28500 35448 29469 35476
rect 28500 35436 28506 35448
rect 29457 35445 29469 35448
rect 29503 35445 29515 35479
rect 29457 35439 29515 35445
rect 30837 35479 30895 35485
rect 30837 35445 30849 35479
rect 30883 35476 30895 35479
rect 31294 35476 31300 35488
rect 30883 35448 31300 35476
rect 30883 35445 30895 35448
rect 30837 35439 30895 35445
rect 31294 35436 31300 35448
rect 31352 35436 31358 35488
rect 31389 35479 31447 35485
rect 31389 35445 31401 35479
rect 31435 35476 31447 35479
rect 32309 35479 32367 35485
rect 32309 35476 32321 35479
rect 31435 35448 32321 35476
rect 31435 35445 31447 35448
rect 31389 35439 31447 35445
rect 32309 35445 32321 35448
rect 32355 35476 32367 35479
rect 32490 35476 32496 35488
rect 32355 35448 32496 35476
rect 32355 35445 32367 35448
rect 32309 35439 32367 35445
rect 32490 35436 32496 35448
rect 32548 35436 32554 35488
rect 33042 35476 33048 35488
rect 33003 35448 33048 35476
rect 33042 35436 33048 35448
rect 33100 35436 33106 35488
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 24394 35272 24400 35284
rect 24355 35244 24400 35272
rect 24394 35232 24400 35244
rect 24452 35232 24458 35284
rect 25314 35232 25320 35284
rect 25372 35272 25378 35284
rect 27157 35275 27215 35281
rect 27157 35272 27169 35275
rect 25372 35244 27169 35272
rect 25372 35232 25378 35244
rect 27157 35241 27169 35244
rect 27203 35241 27215 35275
rect 28626 35272 28632 35284
rect 28587 35244 28632 35272
rect 27157 35235 27215 35241
rect 28626 35232 28632 35244
rect 28684 35232 28690 35284
rect 29641 35275 29699 35281
rect 29641 35241 29653 35275
rect 29687 35272 29699 35275
rect 29822 35272 29828 35284
rect 29687 35244 29828 35272
rect 29687 35241 29699 35244
rect 29641 35235 29699 35241
rect 29822 35232 29828 35244
rect 29880 35272 29886 35284
rect 31662 35272 31668 35284
rect 29880 35244 31668 35272
rect 29880 35232 29886 35244
rect 31662 35232 31668 35244
rect 31720 35232 31726 35284
rect 31941 35275 31999 35281
rect 31941 35241 31953 35275
rect 31987 35272 31999 35275
rect 32122 35272 32128 35284
rect 31987 35244 32128 35272
rect 31987 35241 31999 35244
rect 31941 35235 31999 35241
rect 32122 35232 32128 35244
rect 32180 35232 32186 35284
rect 25869 35207 25927 35213
rect 25869 35173 25881 35207
rect 25915 35204 25927 35207
rect 26418 35204 26424 35216
rect 25915 35176 26424 35204
rect 25915 35173 25927 35176
rect 25869 35167 25927 35173
rect 26418 35164 26424 35176
rect 26476 35164 26482 35216
rect 27798 35204 27804 35216
rect 27759 35176 27804 35204
rect 27798 35164 27804 35176
rect 27856 35164 27862 35216
rect 33042 35204 33048 35216
rect 31726 35176 33048 35204
rect 27341 35139 27399 35145
rect 27341 35136 27353 35139
rect 23676 35108 27353 35136
rect 20162 35068 20168 35080
rect 20123 35040 20168 35068
rect 20162 35028 20168 35040
rect 20220 35028 20226 35080
rect 20349 35071 20407 35077
rect 20349 35037 20361 35071
rect 20395 35068 20407 35071
rect 20438 35068 20444 35080
rect 20395 35040 20444 35068
rect 20395 35037 20407 35040
rect 20349 35031 20407 35037
rect 20438 35028 20444 35040
rect 20496 35028 20502 35080
rect 20806 35068 20812 35080
rect 20767 35040 20812 35068
rect 20806 35028 20812 35040
rect 20864 35028 20870 35080
rect 20990 35068 20996 35080
rect 20951 35040 20996 35068
rect 20990 35028 20996 35040
rect 21048 35028 21054 35080
rect 21818 35028 21824 35080
rect 21876 35068 21882 35080
rect 23676 35077 23704 35108
rect 27341 35105 27353 35108
rect 27387 35136 27399 35139
rect 27614 35136 27620 35148
rect 27387 35108 27620 35136
rect 27387 35105 27399 35108
rect 27341 35099 27399 35105
rect 27614 35096 27620 35108
rect 27672 35096 27678 35148
rect 28810 35096 28816 35148
rect 28868 35136 28874 35148
rect 30926 35136 30932 35148
rect 28868 35108 30932 35136
rect 28868 35096 28874 35108
rect 30926 35096 30932 35108
rect 30984 35096 30990 35148
rect 31726 35136 31754 35176
rect 33042 35164 33048 35176
rect 33100 35164 33106 35216
rect 31312 35108 31754 35136
rect 23661 35071 23719 35077
rect 23661 35068 23673 35071
rect 21876 35040 23673 35068
rect 21876 35028 21882 35040
rect 23661 35037 23673 35040
rect 23707 35037 23719 35071
rect 23842 35068 23848 35080
rect 23803 35040 23848 35068
rect 23661 35031 23719 35037
rect 23842 35028 23848 35040
rect 23900 35028 23906 35080
rect 24026 35028 24032 35080
rect 24084 35068 24090 35080
rect 24394 35068 24400 35080
rect 24084 35040 24400 35068
rect 24084 35028 24090 35040
rect 24394 35028 24400 35040
rect 24452 35068 24458 35080
rect 24555 35071 24613 35077
rect 24555 35068 24567 35071
rect 24452 35040 24567 35068
rect 24452 35028 24458 35040
rect 24555 35037 24567 35040
rect 24601 35037 24613 35071
rect 24555 35031 24613 35037
rect 24662 35071 24720 35077
rect 24662 35037 24674 35071
rect 24708 35037 24720 35071
rect 24662 35031 24720 35037
rect 24765 35071 24823 35077
rect 24765 35037 24777 35071
rect 24811 35037 24823 35071
rect 24765 35031 24823 35037
rect 24857 35071 24915 35077
rect 24857 35037 24869 35071
rect 24903 35068 24915 35071
rect 25498 35068 25504 35080
rect 24903 35040 25504 35068
rect 24903 35037 24915 35040
rect 24857 35031 24915 35037
rect 23750 34960 23756 35012
rect 23808 35000 23814 35012
rect 24688 35000 24716 35031
rect 23808 34972 24716 35000
rect 23808 34960 23814 34972
rect 24780 34944 24808 35031
rect 25498 35028 25504 35040
rect 25556 35028 25562 35080
rect 25682 35028 25688 35080
rect 25740 35068 25746 35080
rect 25777 35071 25835 35077
rect 25777 35068 25789 35071
rect 25740 35040 25789 35068
rect 25740 35028 25746 35040
rect 25777 35037 25789 35040
rect 25823 35037 25835 35071
rect 25777 35031 25835 35037
rect 26053 35071 26111 35077
rect 26053 35037 26065 35071
rect 26099 35037 26111 35071
rect 26053 35031 26111 35037
rect 26068 35000 26096 35031
rect 26142 35028 26148 35080
rect 26200 35068 26206 35080
rect 26237 35071 26295 35077
rect 26237 35068 26249 35071
rect 26200 35040 26249 35068
rect 26200 35028 26206 35040
rect 26237 35037 26249 35040
rect 26283 35037 26295 35071
rect 26237 35031 26295 35037
rect 26418 35028 26424 35080
rect 26476 35068 26482 35080
rect 26513 35071 26571 35077
rect 26513 35068 26525 35071
rect 26476 35040 26525 35068
rect 26476 35028 26482 35040
rect 26513 35037 26525 35040
rect 26559 35037 26571 35071
rect 26513 35031 26571 35037
rect 26602 35028 26608 35080
rect 26660 35068 26666 35080
rect 27065 35071 27123 35077
rect 27065 35068 27077 35071
rect 26660 35040 27077 35068
rect 26660 35028 26666 35040
rect 27065 35037 27077 35040
rect 27111 35037 27123 35071
rect 27065 35031 27123 35037
rect 27801 35071 27859 35077
rect 27801 35037 27813 35071
rect 27847 35068 27859 35071
rect 27890 35068 27896 35080
rect 27847 35040 27896 35068
rect 27847 35037 27859 35040
rect 27801 35031 27859 35037
rect 27890 35028 27896 35040
rect 27948 35028 27954 35080
rect 28074 35068 28080 35080
rect 28035 35040 28080 35068
rect 28074 35028 28080 35040
rect 28132 35028 28138 35080
rect 28534 35068 28540 35080
rect 28495 35040 28540 35068
rect 28534 35028 28540 35040
rect 28592 35028 28598 35080
rect 28721 35071 28779 35077
rect 28721 35037 28733 35071
rect 28767 35037 28779 35071
rect 28721 35031 28779 35037
rect 29917 35071 29975 35077
rect 29917 35037 29929 35071
rect 29963 35068 29975 35071
rect 30282 35068 30288 35080
rect 29963 35040 30288 35068
rect 29963 35037 29975 35040
rect 29917 35031 29975 35037
rect 26326 35000 26332 35012
rect 26068 34972 26332 35000
rect 26326 34960 26332 34972
rect 26384 35000 26390 35012
rect 26970 35000 26976 35012
rect 26384 34972 26976 35000
rect 26384 34960 26390 34972
rect 26970 34960 26976 34972
rect 27028 34960 27034 35012
rect 28442 35000 28448 35012
rect 27908 34972 28448 35000
rect 20254 34932 20260 34944
rect 20215 34904 20260 34932
rect 20254 34892 20260 34904
rect 20312 34892 20318 34944
rect 20346 34892 20352 34944
rect 20404 34932 20410 34944
rect 20901 34935 20959 34941
rect 20901 34932 20913 34935
rect 20404 34904 20913 34932
rect 20404 34892 20410 34904
rect 20901 34901 20913 34904
rect 20947 34901 20959 34935
rect 20901 34895 20959 34901
rect 23845 34935 23903 34941
rect 23845 34901 23857 34935
rect 23891 34932 23903 34935
rect 24670 34932 24676 34944
rect 23891 34904 24676 34932
rect 23891 34901 23903 34904
rect 23845 34895 23903 34901
rect 24670 34892 24676 34904
rect 24728 34892 24734 34944
rect 24762 34892 24768 34944
rect 24820 34892 24826 34944
rect 26418 34892 26424 34944
rect 26476 34932 26482 34944
rect 26786 34932 26792 34944
rect 26476 34904 26792 34932
rect 26476 34892 26482 34904
rect 26786 34892 26792 34904
rect 26844 34892 26850 34944
rect 27341 34935 27399 34941
rect 27341 34901 27353 34935
rect 27387 34932 27399 34935
rect 27908 34932 27936 34972
rect 28442 34960 28448 34972
rect 28500 35000 28506 35012
rect 28736 35000 28764 35031
rect 30282 35028 30288 35040
rect 30340 35028 30346 35080
rect 30374 35028 30380 35080
rect 30432 35028 30438 35080
rect 28500 34972 28764 35000
rect 29641 35003 29699 35009
rect 28500 34960 28506 34972
rect 29641 34969 29653 35003
rect 29687 34969 29699 35003
rect 29641 34963 29699 34969
rect 29825 35003 29883 35009
rect 29825 34969 29837 35003
rect 29871 35000 29883 35003
rect 30392 35000 30420 35028
rect 29871 34972 30420 35000
rect 30837 35003 30895 35009
rect 29871 34969 29883 34972
rect 29825 34963 29883 34969
rect 30837 34969 30849 35003
rect 30883 35000 30895 35003
rect 31312 35000 31340 35108
rect 31570 35068 31576 35080
rect 31531 35040 31576 35068
rect 31570 35028 31576 35040
rect 31628 35028 31634 35080
rect 31662 35028 31668 35080
rect 31720 35068 31726 35080
rect 31757 35071 31815 35077
rect 31757 35068 31769 35071
rect 31720 35040 31769 35068
rect 31720 35028 31726 35040
rect 31757 35037 31769 35040
rect 31803 35037 31815 35071
rect 31757 35031 31815 35037
rect 30883 34972 31340 35000
rect 30883 34969 30895 34972
rect 30837 34963 30895 34969
rect 27387 34904 27936 34932
rect 27387 34901 27399 34904
rect 27341 34895 27399 34901
rect 27982 34892 27988 34944
rect 28040 34932 28046 34944
rect 28040 34904 28085 34932
rect 28040 34892 28046 34904
rect 28166 34892 28172 34944
rect 28224 34932 28230 34944
rect 29656 34932 29684 34963
rect 29730 34932 29736 34944
rect 28224 34904 29736 34932
rect 28224 34892 28230 34904
rect 29730 34892 29736 34904
rect 29788 34932 29794 34944
rect 30190 34932 30196 34944
rect 29788 34904 30196 34932
rect 29788 34892 29794 34904
rect 30190 34892 30196 34904
rect 30248 34892 30254 34944
rect 30377 34935 30435 34941
rect 30377 34901 30389 34935
rect 30423 34932 30435 34935
rect 30466 34932 30472 34944
rect 30423 34904 30472 34932
rect 30423 34901 30435 34904
rect 30377 34895 30435 34901
rect 30466 34892 30472 34904
rect 30524 34892 30530 34944
rect 30745 34935 30803 34941
rect 30745 34901 30757 34935
rect 30791 34932 30803 34935
rect 31386 34932 31392 34944
rect 30791 34904 31392 34932
rect 30791 34901 30803 34904
rect 30745 34895 30803 34901
rect 31386 34892 31392 34904
rect 31444 34892 31450 34944
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 19613 34731 19671 34737
rect 19613 34697 19625 34731
rect 19659 34728 19671 34731
rect 20806 34728 20812 34740
rect 19659 34700 20812 34728
rect 19659 34697 19671 34700
rect 19613 34691 19671 34697
rect 20806 34688 20812 34700
rect 20864 34688 20870 34740
rect 21818 34728 21824 34740
rect 21779 34700 21824 34728
rect 21818 34688 21824 34700
rect 21876 34688 21882 34740
rect 26142 34688 26148 34740
rect 26200 34728 26206 34740
rect 26237 34731 26295 34737
rect 26237 34728 26249 34731
rect 26200 34700 26249 34728
rect 26200 34688 26206 34700
rect 26237 34697 26249 34700
rect 26283 34697 26295 34731
rect 26237 34691 26295 34697
rect 26804 34700 27844 34728
rect 24397 34663 24455 34669
rect 19444 34632 21128 34660
rect 19444 34601 19472 34632
rect 21100 34604 21128 34632
rect 24397 34629 24409 34663
rect 24443 34660 24455 34663
rect 26418 34660 26424 34672
rect 24443 34632 26424 34660
rect 24443 34629 24455 34632
rect 24397 34623 24455 34629
rect 26418 34620 26424 34632
rect 26476 34620 26482 34672
rect 19429 34595 19487 34601
rect 19429 34561 19441 34595
rect 19475 34561 19487 34595
rect 19429 34555 19487 34561
rect 19613 34595 19671 34601
rect 19613 34561 19625 34595
rect 19659 34592 19671 34595
rect 19978 34592 19984 34604
rect 19659 34564 19984 34592
rect 19659 34561 19671 34564
rect 19613 34555 19671 34561
rect 19978 34552 19984 34564
rect 20036 34552 20042 34604
rect 20254 34592 20260 34604
rect 20215 34564 20260 34592
rect 20254 34552 20260 34564
rect 20312 34552 20318 34604
rect 21082 34592 21088 34604
rect 20995 34564 21088 34592
rect 21082 34552 21088 34564
rect 21140 34552 21146 34604
rect 21177 34595 21235 34601
rect 21177 34561 21189 34595
rect 21223 34592 21235 34595
rect 22189 34595 22247 34601
rect 22189 34592 22201 34595
rect 21223 34564 22201 34592
rect 21223 34561 21235 34564
rect 21177 34555 21235 34561
rect 22189 34561 22201 34564
rect 22235 34561 22247 34595
rect 22189 34555 22247 34561
rect 23658 34552 23664 34604
rect 23716 34552 23722 34604
rect 24670 34552 24676 34604
rect 24728 34592 24734 34604
rect 24854 34592 24860 34604
rect 24728 34564 24860 34592
rect 24728 34552 24734 34564
rect 24854 34552 24860 34564
rect 24912 34552 24918 34604
rect 25314 34552 25320 34604
rect 25372 34592 25378 34604
rect 25866 34592 25872 34604
rect 25372 34564 25872 34592
rect 25372 34552 25378 34564
rect 25866 34552 25872 34564
rect 25924 34592 25930 34604
rect 26145 34595 26203 34601
rect 26145 34592 26157 34595
rect 25924 34564 26157 34592
rect 25924 34552 25930 34564
rect 26145 34561 26157 34564
rect 26191 34561 26203 34595
rect 26145 34555 26203 34561
rect 26329 34595 26387 34601
rect 26329 34561 26341 34595
rect 26375 34592 26387 34595
rect 26510 34592 26516 34604
rect 26375 34564 26516 34592
rect 26375 34561 26387 34564
rect 26329 34555 26387 34561
rect 26510 34552 26516 34564
rect 26568 34552 26574 34604
rect 20346 34524 20352 34536
rect 20307 34496 20352 34524
rect 20346 34484 20352 34496
rect 20404 34484 20410 34536
rect 22281 34527 22339 34533
rect 22281 34524 22293 34527
rect 21376 34496 22293 34524
rect 20625 34459 20683 34465
rect 20625 34425 20637 34459
rect 20671 34456 20683 34459
rect 21376 34456 21404 34496
rect 22281 34493 22293 34496
rect 22327 34493 22339 34527
rect 22281 34487 22339 34493
rect 22465 34527 22523 34533
rect 22465 34493 22477 34527
rect 22511 34493 22523 34527
rect 23566 34524 23572 34536
rect 23527 34496 23572 34524
rect 22465 34487 22523 34493
rect 20671 34428 21404 34456
rect 22480 34456 22508 34487
rect 23566 34484 23572 34496
rect 23624 34484 23630 34536
rect 23750 34484 23756 34536
rect 23808 34524 23814 34536
rect 25133 34527 25191 34533
rect 25133 34524 25145 34527
rect 23808 34496 25145 34524
rect 23808 34484 23814 34496
rect 24044 34468 24072 34496
rect 25133 34493 25145 34496
rect 25179 34524 25191 34527
rect 26804 34524 26832 34700
rect 27706 34660 27712 34672
rect 27172 34632 27712 34660
rect 26878 34552 26884 34604
rect 26936 34592 26942 34604
rect 27172 34601 27200 34632
rect 27706 34620 27712 34632
rect 27764 34620 27770 34672
rect 27816 34660 27844 34700
rect 27890 34688 27896 34740
rect 27948 34728 27954 34740
rect 30561 34731 30619 34737
rect 27948 34700 28580 34728
rect 27948 34688 27954 34700
rect 28552 34672 28580 34700
rect 30561 34697 30573 34731
rect 30607 34728 30619 34731
rect 31386 34728 31392 34740
rect 30607 34700 31248 34728
rect 31347 34700 31392 34728
rect 30607 34697 30619 34700
rect 30561 34691 30619 34697
rect 27982 34660 27988 34672
rect 27816 34632 27988 34660
rect 27982 34620 27988 34632
rect 28040 34660 28046 34672
rect 28445 34663 28503 34669
rect 28445 34660 28457 34663
rect 28040 34632 28457 34660
rect 28040 34620 28046 34632
rect 28445 34629 28457 34632
rect 28491 34629 28503 34663
rect 28445 34623 28503 34629
rect 28534 34620 28540 34672
rect 28592 34660 28598 34672
rect 28645 34663 28703 34669
rect 28645 34660 28657 34663
rect 28592 34632 28657 34660
rect 28592 34620 28598 34632
rect 28645 34629 28657 34632
rect 28691 34629 28703 34663
rect 30190 34660 30196 34672
rect 30151 34632 30196 34660
rect 28645 34623 28703 34629
rect 30190 34620 30196 34632
rect 30248 34620 30254 34672
rect 30282 34620 30288 34672
rect 30340 34660 30346 34672
rect 30393 34663 30451 34669
rect 30393 34660 30405 34663
rect 30340 34632 30405 34660
rect 30340 34620 30346 34632
rect 30393 34629 30405 34632
rect 30439 34660 30451 34663
rect 31220 34660 31248 34700
rect 31386 34688 31392 34700
rect 31444 34688 31450 34740
rect 31570 34660 31576 34672
rect 30439 34632 31156 34660
rect 31220 34632 31576 34660
rect 30439 34629 30451 34632
rect 30393 34623 30451 34629
rect 26973 34595 27031 34601
rect 26973 34592 26985 34595
rect 26936 34564 26985 34592
rect 26936 34552 26942 34564
rect 26973 34561 26985 34564
rect 27019 34561 27031 34595
rect 26973 34555 27031 34561
rect 27157 34595 27215 34601
rect 27157 34561 27169 34595
rect 27203 34561 27215 34595
rect 27614 34592 27620 34604
rect 27575 34564 27620 34592
rect 27157 34555 27215 34561
rect 27614 34552 27620 34564
rect 27672 34552 27678 34604
rect 27801 34595 27859 34601
rect 27801 34561 27813 34595
rect 27847 34592 27859 34595
rect 28166 34592 28172 34604
rect 27847 34564 28172 34592
rect 27847 34561 27859 34564
rect 27801 34555 27859 34561
rect 28166 34552 28172 34564
rect 28224 34552 28230 34604
rect 29270 34592 29276 34604
rect 29231 34564 29276 34592
rect 29270 34552 29276 34564
rect 29328 34552 29334 34604
rect 29454 34592 29460 34604
rect 29415 34564 29460 34592
rect 29454 34552 29460 34564
rect 29512 34552 29518 34604
rect 31018 34592 31024 34604
rect 30979 34564 31024 34592
rect 31018 34552 31024 34564
rect 31076 34552 31082 34604
rect 31128 34592 31156 34632
rect 31570 34620 31576 34632
rect 31628 34620 31634 34672
rect 34606 34660 34612 34672
rect 32048 34632 34612 34660
rect 31205 34595 31263 34601
rect 31205 34592 31217 34595
rect 31128 34564 31217 34592
rect 31205 34561 31217 34564
rect 31251 34561 31263 34595
rect 31205 34555 31263 34561
rect 25179 34496 26832 34524
rect 27065 34527 27123 34533
rect 25179 34493 25191 34496
rect 25133 34487 25191 34493
rect 27065 34493 27077 34527
rect 27111 34524 27123 34527
rect 32048 34524 32076 34632
rect 34606 34620 34612 34632
rect 34664 34620 34670 34672
rect 32125 34595 32183 34601
rect 32125 34561 32137 34595
rect 32171 34592 32183 34595
rect 32214 34592 32220 34604
rect 32171 34564 32220 34592
rect 32171 34561 32183 34564
rect 32125 34555 32183 34561
rect 32214 34552 32220 34564
rect 32272 34552 32278 34604
rect 37829 34595 37887 34601
rect 37829 34561 37841 34595
rect 37875 34592 37887 34595
rect 38194 34592 38200 34604
rect 37875 34564 38200 34592
rect 37875 34561 37887 34564
rect 37829 34555 37887 34561
rect 38194 34552 38200 34564
rect 38252 34552 38258 34604
rect 32398 34524 32404 34536
rect 27111 34496 32076 34524
rect 32359 34496 32404 34524
rect 27111 34493 27123 34496
rect 27065 34487 27123 34493
rect 32398 34484 32404 34496
rect 32456 34484 32462 34536
rect 22830 34456 22836 34468
rect 22480 34428 22836 34456
rect 20671 34425 20683 34428
rect 20625 34419 20683 34425
rect 22830 34416 22836 34428
rect 22888 34416 22894 34468
rect 24026 34416 24032 34468
rect 24084 34416 24090 34468
rect 27985 34391 28043 34397
rect 27985 34357 27997 34391
rect 28031 34388 28043 34391
rect 28074 34388 28080 34400
rect 28031 34360 28080 34388
rect 28031 34357 28043 34360
rect 27985 34351 28043 34357
rect 28074 34348 28080 34360
rect 28132 34388 28138 34400
rect 28626 34388 28632 34400
rect 28132 34360 28632 34388
rect 28132 34348 28138 34360
rect 28626 34348 28632 34360
rect 28684 34348 28690 34400
rect 28810 34388 28816 34400
rect 28771 34360 28816 34388
rect 28810 34348 28816 34360
rect 28868 34348 28874 34400
rect 29273 34391 29331 34397
rect 29273 34357 29285 34391
rect 29319 34388 29331 34391
rect 29822 34388 29828 34400
rect 29319 34360 29828 34388
rect 29319 34357 29331 34360
rect 29273 34351 29331 34357
rect 29822 34348 29828 34360
rect 29880 34348 29886 34400
rect 30374 34388 30380 34400
rect 30335 34360 30380 34388
rect 30374 34348 30380 34360
rect 30432 34388 30438 34400
rect 31018 34388 31024 34400
rect 30432 34360 31024 34388
rect 30432 34348 30438 34360
rect 31018 34348 31024 34360
rect 31076 34348 31082 34400
rect 31386 34348 31392 34400
rect 31444 34388 31450 34400
rect 31754 34388 31760 34400
rect 31444 34360 31760 34388
rect 31444 34348 31450 34360
rect 31754 34348 31760 34360
rect 31812 34388 31818 34400
rect 32217 34391 32275 34397
rect 32217 34388 32229 34391
rect 31812 34360 32229 34388
rect 31812 34348 31818 34360
rect 32217 34357 32229 34360
rect 32263 34357 32275 34391
rect 32217 34351 32275 34357
rect 32306 34348 32312 34400
rect 32364 34388 32370 34400
rect 38010 34388 38016 34400
rect 32364 34360 32409 34388
rect 37971 34360 38016 34388
rect 32364 34348 32370 34360
rect 38010 34348 38016 34360
rect 38068 34348 38074 34400
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 19797 34187 19855 34193
rect 19797 34153 19809 34187
rect 19843 34184 19855 34187
rect 19843 34156 20116 34184
rect 19843 34153 19855 34156
rect 19797 34147 19855 34153
rect 20088 34128 20116 34156
rect 21082 34144 21088 34196
rect 21140 34184 21146 34196
rect 21637 34187 21695 34193
rect 21637 34184 21649 34187
rect 21140 34156 21649 34184
rect 21140 34144 21146 34156
rect 21637 34153 21649 34156
rect 21683 34153 21695 34187
rect 21637 34147 21695 34153
rect 25590 34144 25596 34196
rect 25648 34184 25654 34196
rect 28169 34187 28227 34193
rect 28169 34184 28181 34187
rect 25648 34156 28181 34184
rect 25648 34144 25654 34156
rect 28169 34153 28181 34156
rect 28215 34153 28227 34187
rect 28169 34147 28227 34153
rect 19981 34119 20039 34125
rect 19981 34085 19993 34119
rect 20027 34085 20039 34119
rect 19981 34079 20039 34085
rect 19996 34048 20024 34079
rect 20070 34076 20076 34128
rect 20128 34116 20134 34128
rect 26145 34119 26203 34125
rect 20128 34088 21496 34116
rect 20128 34076 20134 34088
rect 20625 34051 20683 34057
rect 20625 34048 20637 34051
rect 19996 34020 20637 34048
rect 20625 34017 20637 34020
rect 20671 34048 20683 34051
rect 20990 34048 20996 34060
rect 20671 34020 20996 34048
rect 20671 34017 20683 34020
rect 20625 34011 20683 34017
rect 20990 34008 20996 34020
rect 21048 34008 21054 34060
rect 19242 33940 19248 33992
rect 19300 33980 19306 33992
rect 19613 33983 19671 33989
rect 19613 33980 19625 33983
rect 19300 33952 19625 33980
rect 19300 33940 19306 33952
rect 19613 33949 19625 33952
rect 19659 33949 19671 33983
rect 19613 33943 19671 33949
rect 19797 33983 19855 33989
rect 19797 33949 19809 33983
rect 19843 33980 19855 33983
rect 19978 33980 19984 33992
rect 19843 33952 19984 33980
rect 19843 33949 19855 33952
rect 19797 33943 19855 33949
rect 19628 33912 19656 33943
rect 19978 33940 19984 33952
rect 20036 33940 20042 33992
rect 20254 33940 20260 33992
rect 20312 33980 20318 33992
rect 20441 33983 20499 33989
rect 20441 33980 20453 33983
rect 20312 33952 20453 33980
rect 20312 33940 20318 33952
rect 20441 33949 20453 33952
rect 20487 33949 20499 33983
rect 20806 33980 20812 33992
rect 20767 33952 20812 33980
rect 20441 33943 20499 33949
rect 20806 33940 20812 33952
rect 20864 33940 20870 33992
rect 21468 33989 21496 34088
rect 26145 34085 26157 34119
rect 26191 34085 26203 34119
rect 28184 34116 28212 34147
rect 28442 34144 28448 34196
rect 28500 34184 28506 34196
rect 28629 34187 28687 34193
rect 28629 34184 28641 34187
rect 28500 34156 28641 34184
rect 28500 34144 28506 34156
rect 28629 34153 28641 34156
rect 28675 34153 28687 34187
rect 29638 34184 29644 34196
rect 28629 34147 28687 34153
rect 28828 34156 29644 34184
rect 28828 34116 28856 34156
rect 29638 34144 29644 34156
rect 29696 34144 29702 34196
rect 29825 34187 29883 34193
rect 29825 34153 29837 34187
rect 29871 34184 29883 34187
rect 29914 34184 29920 34196
rect 29871 34156 29920 34184
rect 29871 34153 29883 34156
rect 29825 34147 29883 34153
rect 29840 34116 29868 34147
rect 29914 34144 29920 34156
rect 29972 34144 29978 34196
rect 30009 34187 30067 34193
rect 30009 34153 30021 34187
rect 30055 34184 30067 34187
rect 30282 34184 30288 34196
rect 30055 34156 30288 34184
rect 30055 34153 30067 34156
rect 30009 34147 30067 34153
rect 30282 34144 30288 34156
rect 30340 34144 30346 34196
rect 31297 34187 31355 34193
rect 31297 34153 31309 34187
rect 31343 34184 31355 34187
rect 31386 34184 31392 34196
rect 31343 34156 31392 34184
rect 31343 34153 31355 34156
rect 31297 34147 31355 34153
rect 31386 34144 31392 34156
rect 31444 34144 31450 34196
rect 28184 34088 28856 34116
rect 28920 34088 29868 34116
rect 26145 34079 26203 34085
rect 23566 34008 23572 34060
rect 23624 34048 23630 34060
rect 23845 34051 23903 34057
rect 23845 34048 23857 34051
rect 23624 34020 23857 34048
rect 23624 34008 23630 34020
rect 23845 34017 23857 34020
rect 23891 34048 23903 34051
rect 24118 34048 24124 34060
rect 23891 34020 24124 34048
rect 23891 34017 23903 34020
rect 23845 34011 23903 34017
rect 24118 34008 24124 34020
rect 24176 34048 24182 34060
rect 24762 34048 24768 34060
rect 24176 34020 24768 34048
rect 24176 34008 24182 34020
rect 24762 34008 24768 34020
rect 24820 34048 24826 34060
rect 25498 34048 25504 34060
rect 24820 34020 25176 34048
rect 25459 34020 25504 34048
rect 24820 34008 24826 34020
rect 21453 33983 21511 33989
rect 21453 33949 21465 33983
rect 21499 33949 21511 33983
rect 23474 33980 23480 33992
rect 23435 33952 23480 33980
rect 21453 33943 21511 33949
rect 23474 33940 23480 33952
rect 23532 33940 23538 33992
rect 23750 33980 23756 33992
rect 23711 33952 23756 33980
rect 23750 33940 23756 33952
rect 23808 33940 23814 33992
rect 24673 33983 24731 33989
rect 24673 33949 24685 33983
rect 24719 33949 24731 33983
rect 24854 33980 24860 33992
rect 24815 33952 24860 33980
rect 24673 33943 24731 33949
rect 21269 33915 21327 33921
rect 21269 33912 21281 33915
rect 19628 33884 21281 33912
rect 21269 33881 21281 33884
rect 21315 33881 21327 33915
rect 21269 33875 21327 33881
rect 23934 33872 23940 33924
rect 23992 33912 23998 33924
rect 24394 33912 24400 33924
rect 23992 33884 24400 33912
rect 23992 33872 23998 33884
rect 24394 33872 24400 33884
rect 24452 33912 24458 33924
rect 24688 33912 24716 33943
rect 24854 33940 24860 33952
rect 24912 33940 24918 33992
rect 25148 33989 25176 34020
rect 25498 34008 25504 34020
rect 25556 34008 25562 34060
rect 26160 34048 26188 34079
rect 26697 34051 26755 34057
rect 26697 34048 26709 34051
rect 26160 34020 26709 34048
rect 26697 34017 26709 34020
rect 26743 34048 26755 34051
rect 28353 34051 28411 34057
rect 26743 34020 28304 34048
rect 26743 34017 26755 34020
rect 26697 34011 26755 34017
rect 25133 33983 25191 33989
rect 25133 33949 25145 33983
rect 25179 33949 25191 33983
rect 25958 33980 25964 33992
rect 25919 33952 25964 33980
rect 25133 33943 25191 33949
rect 25958 33940 25964 33952
rect 26016 33940 26022 33992
rect 26510 33940 26516 33992
rect 26568 33980 26574 33992
rect 26973 33983 27031 33989
rect 26973 33980 26985 33983
rect 26568 33952 26985 33980
rect 26568 33940 26574 33952
rect 26973 33949 26985 33952
rect 27019 33980 27031 33983
rect 27430 33980 27436 33992
rect 27019 33952 27436 33980
rect 27019 33949 27031 33952
rect 26973 33943 27031 33949
rect 27430 33940 27436 33952
rect 27488 33940 27494 33992
rect 27798 33940 27804 33992
rect 27856 33980 27862 33992
rect 28169 33983 28227 33989
rect 28169 33980 28181 33983
rect 27856 33952 28181 33980
rect 27856 33940 27862 33952
rect 28169 33949 28181 33952
rect 28215 33949 28227 33983
rect 28276 33980 28304 34020
rect 28353 34017 28365 34051
rect 28399 34048 28411 34051
rect 28810 34048 28816 34060
rect 28399 34020 28816 34048
rect 28399 34017 28411 34020
rect 28353 34011 28411 34017
rect 28810 34008 28816 34020
rect 28868 34008 28874 34060
rect 28445 33983 28503 33989
rect 28445 33980 28457 33983
rect 28276 33952 28457 33980
rect 28169 33943 28227 33949
rect 28445 33949 28457 33952
rect 28491 33980 28503 33983
rect 28920 33980 28948 34088
rect 31662 34076 31668 34128
rect 31720 34116 31726 34128
rect 31938 34116 31944 34128
rect 31720 34088 31944 34116
rect 31720 34076 31726 34088
rect 31938 34076 31944 34088
rect 31996 34076 32002 34128
rect 32953 34119 33011 34125
rect 32953 34116 32965 34119
rect 32416 34088 32965 34116
rect 32416 34060 32444 34088
rect 32953 34085 32965 34088
rect 32999 34085 33011 34119
rect 32953 34079 33011 34085
rect 29638 34048 29644 34060
rect 29599 34020 29644 34048
rect 29638 34008 29644 34020
rect 29696 34008 29702 34060
rect 32398 34048 32404 34060
rect 31128 34020 32404 34048
rect 29822 33980 29828 33992
rect 28491 33952 28948 33980
rect 29783 33952 29828 33980
rect 28491 33949 28503 33952
rect 28445 33943 28503 33949
rect 29822 33940 29828 33952
rect 29880 33940 29886 33992
rect 30469 33983 30527 33989
rect 30469 33949 30481 33983
rect 30515 33949 30527 33983
rect 30469 33943 30527 33949
rect 30653 33983 30711 33989
rect 30653 33949 30665 33983
rect 30699 33980 30711 33983
rect 30742 33980 30748 33992
rect 30699 33952 30748 33980
rect 30699 33949 30711 33952
rect 30653 33943 30711 33949
rect 28718 33912 28724 33924
rect 24452 33884 28724 33912
rect 24452 33872 24458 33884
rect 28718 33872 28724 33884
rect 28776 33872 28782 33924
rect 29549 33915 29607 33921
rect 29549 33881 29561 33915
rect 29595 33912 29607 33915
rect 30282 33912 30288 33924
rect 29595 33884 30288 33912
rect 29595 33881 29607 33884
rect 29549 33875 29607 33881
rect 30282 33872 30288 33884
rect 30340 33872 30346 33924
rect 30484 33912 30512 33943
rect 30742 33940 30748 33952
rect 30800 33940 30806 33992
rect 31128 33989 31156 34020
rect 32398 34008 32404 34020
rect 32456 34008 32462 34060
rect 33042 34048 33048 34060
rect 33003 34020 33048 34048
rect 33042 34008 33048 34020
rect 33100 34008 33106 34060
rect 31113 33983 31171 33989
rect 31113 33949 31125 33983
rect 31159 33949 31171 33983
rect 31113 33943 31171 33949
rect 31297 33983 31355 33989
rect 31297 33949 31309 33983
rect 31343 33980 31355 33983
rect 31938 33980 31944 33992
rect 31343 33952 31754 33980
rect 31899 33952 31944 33980
rect 31343 33949 31355 33952
rect 31297 33943 31355 33949
rect 31726 33912 31754 33952
rect 31938 33940 31944 33952
rect 31996 33940 32002 33992
rect 32125 33983 32183 33989
rect 32125 33949 32137 33983
rect 32171 33980 32183 33983
rect 32766 33980 32772 33992
rect 32171 33952 32444 33980
rect 32727 33952 32772 33980
rect 32171 33949 32183 33952
rect 32125 33943 32183 33949
rect 32214 33912 32220 33924
rect 30484 33884 31616 33912
rect 31726 33884 32220 33912
rect 20346 33804 20352 33856
rect 20404 33844 20410 33856
rect 20533 33847 20591 33853
rect 20533 33844 20545 33847
rect 20404 33816 20545 33844
rect 20404 33804 20410 33816
rect 20533 33813 20545 33816
rect 20579 33813 20591 33847
rect 20714 33844 20720 33856
rect 20675 33816 20720 33844
rect 20533 33807 20591 33813
rect 20714 33804 20720 33816
rect 20772 33804 20778 33856
rect 30190 33804 30196 33856
rect 30248 33844 30254 33856
rect 30484 33844 30512 33884
rect 30248 33816 30512 33844
rect 30561 33847 30619 33853
rect 30248 33804 30254 33816
rect 30561 33813 30573 33847
rect 30607 33844 30619 33847
rect 30834 33844 30840 33856
rect 30607 33816 30840 33844
rect 30607 33813 30619 33816
rect 30561 33807 30619 33813
rect 30834 33804 30840 33816
rect 30892 33804 30898 33856
rect 31202 33804 31208 33856
rect 31260 33844 31266 33856
rect 31481 33847 31539 33853
rect 31481 33844 31493 33847
rect 31260 33816 31493 33844
rect 31260 33804 31266 33816
rect 31481 33813 31493 33816
rect 31527 33813 31539 33847
rect 31588 33844 31616 33884
rect 32214 33872 32220 33884
rect 32272 33912 32278 33924
rect 32309 33915 32367 33921
rect 32309 33912 32321 33915
rect 32272 33884 32321 33912
rect 32272 33872 32278 33884
rect 32309 33881 32321 33884
rect 32355 33881 32367 33915
rect 32416 33912 32444 33952
rect 32766 33940 32772 33952
rect 32824 33940 32830 33992
rect 32861 33983 32919 33989
rect 32861 33949 32873 33983
rect 32907 33980 32919 33983
rect 33870 33980 33876 33992
rect 32907 33952 33876 33980
rect 32907 33949 32919 33952
rect 32861 33943 32919 33949
rect 33870 33940 33876 33952
rect 33928 33940 33934 33992
rect 32674 33912 32680 33924
rect 32416 33884 32680 33912
rect 32309 33875 32367 33881
rect 32674 33872 32680 33884
rect 32732 33872 32738 33924
rect 31662 33844 31668 33856
rect 31588 33816 31668 33844
rect 31481 33807 31539 33813
rect 31662 33804 31668 33816
rect 31720 33804 31726 33856
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 20990 33640 20996 33652
rect 20456 33612 20996 33640
rect 20456 33581 20484 33612
rect 20990 33600 20996 33612
rect 21048 33600 21054 33652
rect 24949 33643 25007 33649
rect 24949 33609 24961 33643
rect 24995 33640 25007 33643
rect 25958 33640 25964 33652
rect 24995 33612 25964 33640
rect 24995 33609 25007 33612
rect 24949 33603 25007 33609
rect 20441 33575 20499 33581
rect 20441 33541 20453 33575
rect 20487 33541 20499 33575
rect 20806 33572 20812 33584
rect 20441 33535 20499 33541
rect 20640 33544 20812 33572
rect 19337 33507 19395 33513
rect 19337 33473 19349 33507
rect 19383 33473 19395 33507
rect 19337 33467 19395 33473
rect 19352 33436 19380 33467
rect 19426 33464 19432 33516
rect 19484 33504 19490 33516
rect 19613 33507 19671 33513
rect 19613 33504 19625 33507
rect 19484 33476 19625 33504
rect 19484 33464 19490 33476
rect 19613 33473 19625 33476
rect 19659 33504 19671 33507
rect 20070 33504 20076 33516
rect 19659 33476 20076 33504
rect 19659 33473 19671 33476
rect 19613 33467 19671 33473
rect 20070 33464 20076 33476
rect 20128 33464 20134 33516
rect 20254 33504 20260 33516
rect 20215 33476 20260 33504
rect 20254 33464 20260 33476
rect 20312 33464 20318 33516
rect 20346 33464 20352 33516
rect 20404 33504 20410 33516
rect 20640 33513 20668 33544
rect 20806 33532 20812 33544
rect 20864 33532 20870 33584
rect 24118 33572 24124 33584
rect 24079 33544 24124 33572
rect 24118 33532 24124 33544
rect 24176 33532 24182 33584
rect 24964 33572 24992 33603
rect 25958 33600 25964 33612
rect 26016 33600 26022 33652
rect 26970 33640 26976 33652
rect 26931 33612 26976 33640
rect 26970 33600 26976 33612
rect 27028 33600 27034 33652
rect 30282 33640 30288 33652
rect 30243 33612 30288 33640
rect 30282 33600 30288 33612
rect 30340 33600 30346 33652
rect 29270 33572 29276 33584
rect 24412 33544 24992 33572
rect 28460 33544 29276 33572
rect 20625 33507 20683 33513
rect 20404 33476 20449 33504
rect 20404 33464 20410 33476
rect 20625 33473 20637 33507
rect 20671 33473 20683 33507
rect 20625 33467 20683 33473
rect 20717 33507 20775 33513
rect 20717 33473 20729 33507
rect 20763 33473 20775 33507
rect 22186 33504 22192 33516
rect 22147 33476 22192 33504
rect 20717 33467 20775 33473
rect 19978 33436 19984 33448
rect 19352 33408 19984 33436
rect 19978 33396 19984 33408
rect 20036 33436 20042 33448
rect 20438 33436 20444 33448
rect 20036 33408 20444 33436
rect 20036 33396 20042 33408
rect 20438 33396 20444 33408
rect 20496 33396 20502 33448
rect 19153 33371 19211 33377
rect 19153 33337 19165 33371
rect 19199 33368 19211 33371
rect 20640 33368 20668 33467
rect 20732 33436 20760 33467
rect 22186 33464 22192 33476
rect 22244 33464 22250 33516
rect 23934 33504 23940 33516
rect 23895 33476 23940 33504
rect 23934 33464 23940 33476
rect 23992 33464 23998 33516
rect 24026 33464 24032 33516
rect 24084 33504 24090 33516
rect 24412 33513 24440 33544
rect 28460 33516 28488 33544
rect 29270 33532 29276 33544
rect 29328 33572 29334 33584
rect 31202 33572 31208 33584
rect 29328 33544 30144 33572
rect 31163 33544 31208 33572
rect 29328 33532 29334 33544
rect 24305 33507 24363 33513
rect 24084 33476 24129 33504
rect 24084 33464 24090 33476
rect 24305 33473 24317 33507
rect 24351 33473 24363 33507
rect 24305 33467 24363 33473
rect 24397 33507 24455 33513
rect 24397 33473 24409 33507
rect 24443 33473 24455 33507
rect 24854 33504 24860 33516
rect 24815 33476 24860 33504
rect 24397 33467 24455 33473
rect 20806 33436 20812 33448
rect 20732 33408 20812 33436
rect 20806 33396 20812 33408
rect 20864 33396 20870 33448
rect 22278 33436 22284 33448
rect 22239 33408 22284 33436
rect 22278 33396 22284 33408
rect 22336 33396 22342 33448
rect 22465 33439 22523 33445
rect 22465 33405 22477 33439
rect 22511 33436 22523 33439
rect 22830 33436 22836 33448
rect 22511 33408 22836 33436
rect 22511 33405 22523 33408
rect 22465 33399 22523 33405
rect 22830 33396 22836 33408
rect 22888 33396 22894 33448
rect 23474 33396 23480 33448
rect 23532 33436 23538 33448
rect 24320 33436 24348 33467
rect 24854 33464 24860 33476
rect 24912 33464 24918 33516
rect 25041 33507 25099 33513
rect 25041 33473 25053 33507
rect 25087 33504 25099 33507
rect 25774 33504 25780 33516
rect 25087 33476 25780 33504
rect 25087 33473 25099 33476
rect 25041 33467 25099 33473
rect 25774 33464 25780 33476
rect 25832 33464 25838 33516
rect 25866 33464 25872 33516
rect 25924 33504 25930 33516
rect 25924 33476 25969 33504
rect 25924 33464 25930 33476
rect 26050 33464 26056 33516
rect 26108 33504 26114 33516
rect 27157 33507 27215 33513
rect 27157 33504 27169 33507
rect 26108 33476 27169 33504
rect 26108 33464 26114 33476
rect 27157 33473 27169 33476
rect 27203 33473 27215 33507
rect 27430 33504 27436 33516
rect 27391 33476 27436 33504
rect 27157 33467 27215 33473
rect 27430 33464 27436 33476
rect 27488 33464 27494 33516
rect 28442 33504 28448 33516
rect 28403 33476 28448 33504
rect 28442 33464 28448 33476
rect 28500 33464 28506 33516
rect 28626 33464 28632 33516
rect 28684 33504 28690 33516
rect 28721 33507 28779 33513
rect 28721 33504 28733 33507
rect 28684 33476 28733 33504
rect 28684 33464 28690 33476
rect 28721 33473 28733 33476
rect 28767 33473 28779 33507
rect 29086 33504 29092 33516
rect 29047 33476 29092 33504
rect 28721 33467 28779 33473
rect 29086 33464 29092 33476
rect 29144 33464 29150 33516
rect 29454 33464 29460 33516
rect 29512 33504 29518 33516
rect 30116 33513 30144 33544
rect 31202 33532 31208 33544
rect 31260 33532 31266 33584
rect 31662 33572 31668 33584
rect 31312 33544 31668 33572
rect 31312 33516 31340 33544
rect 31662 33532 31668 33544
rect 31720 33532 31726 33584
rect 32766 33532 32772 33584
rect 32824 33572 32830 33584
rect 32824 33544 34008 33572
rect 32824 33532 32830 33544
rect 29917 33507 29975 33513
rect 29917 33504 29929 33507
rect 29512 33476 29929 33504
rect 29512 33464 29518 33476
rect 29917 33473 29929 33476
rect 29963 33473 29975 33507
rect 29917 33467 29975 33473
rect 30101 33507 30159 33513
rect 30101 33473 30113 33507
rect 30147 33473 30159 33507
rect 30101 33467 30159 33473
rect 30929 33507 30987 33513
rect 30929 33473 30941 33507
rect 30975 33473 30987 33507
rect 30929 33467 30987 33473
rect 31077 33507 31135 33513
rect 31077 33473 31089 33507
rect 31123 33504 31135 33507
rect 31294 33504 31300 33516
rect 31123 33473 31156 33504
rect 31255 33476 31300 33504
rect 31077 33467 31156 33473
rect 24670 33436 24676 33448
rect 23532 33408 24676 33436
rect 23532 33396 23538 33408
rect 24670 33396 24676 33408
rect 24728 33436 24734 33448
rect 25498 33436 25504 33448
rect 24728 33408 25504 33436
rect 24728 33396 24734 33408
rect 25498 33396 25504 33408
rect 25556 33396 25562 33448
rect 25590 33396 25596 33448
rect 25648 33436 25654 33448
rect 25884 33436 25912 33464
rect 27341 33439 27399 33445
rect 27341 33436 27353 33439
rect 25648 33408 25693 33436
rect 25884 33408 27353 33436
rect 25648 33396 25654 33408
rect 27341 33405 27353 33408
rect 27387 33405 27399 33439
rect 27341 33399 27399 33405
rect 28169 33439 28227 33445
rect 28169 33405 28181 33439
rect 28215 33436 28227 33439
rect 28994 33436 29000 33448
rect 28215 33408 29000 33436
rect 28215 33405 28227 33408
rect 28169 33399 28227 33405
rect 28994 33396 29000 33408
rect 29052 33436 29058 33448
rect 29472 33436 29500 33464
rect 29052 33408 29500 33436
rect 29052 33396 29058 33408
rect 19199 33340 20668 33368
rect 19199 33337 19211 33340
rect 19153 33331 19211 33337
rect 24854 33328 24860 33380
rect 24912 33368 24918 33380
rect 25038 33368 25044 33380
rect 24912 33340 25044 33368
rect 24912 33328 24918 33340
rect 25038 33328 25044 33340
rect 25096 33328 25102 33380
rect 28718 33368 28724 33380
rect 28679 33340 28724 33368
rect 28718 33328 28724 33340
rect 28776 33328 28782 33380
rect 30944 33368 30972 33467
rect 31128 33436 31156 33467
rect 31294 33464 31300 33476
rect 31352 33464 31358 33516
rect 31386 33464 31392 33516
rect 31444 33513 31450 33516
rect 31444 33507 31471 33513
rect 31459 33473 31471 33507
rect 31444 33467 31471 33473
rect 31444 33464 31450 33467
rect 31938 33464 31944 33516
rect 31996 33504 32002 33516
rect 32493 33507 32551 33513
rect 32493 33504 32505 33507
rect 31996 33476 32505 33504
rect 31996 33464 32002 33476
rect 32493 33473 32505 33476
rect 32539 33504 32551 33507
rect 32858 33504 32864 33516
rect 32539 33476 32864 33504
rect 32539 33473 32551 33476
rect 32493 33467 32551 33473
rect 32858 33464 32864 33476
rect 32916 33464 32922 33516
rect 33980 33513 34008 33544
rect 33965 33507 34023 33513
rect 33965 33473 33977 33507
rect 34011 33473 34023 33507
rect 33965 33467 34023 33473
rect 32306 33436 32312 33448
rect 31128 33408 32312 33436
rect 32306 33396 32312 33408
rect 32364 33396 32370 33448
rect 32769 33439 32827 33445
rect 32769 33405 32781 33439
rect 32815 33405 32827 33439
rect 33870 33436 33876 33448
rect 33831 33408 33876 33436
rect 32769 33399 32827 33405
rect 30944 33340 31754 33368
rect 18322 33260 18328 33312
rect 18380 33300 18386 33312
rect 19242 33300 19248 33312
rect 18380 33272 19248 33300
rect 18380 33260 18386 33272
rect 19242 33260 19248 33272
rect 19300 33300 19306 33312
rect 19521 33303 19579 33309
rect 19521 33300 19533 33303
rect 19300 33272 19533 33300
rect 19300 33260 19306 33272
rect 19521 33269 19533 33272
rect 19567 33269 19579 33303
rect 19521 33263 19579 33269
rect 20073 33303 20131 33309
rect 20073 33269 20085 33303
rect 20119 33300 20131 33303
rect 21082 33300 21088 33312
rect 20119 33272 21088 33300
rect 20119 33269 20131 33272
rect 20073 33263 20131 33269
rect 21082 33260 21088 33272
rect 21140 33260 21146 33312
rect 21821 33303 21879 33309
rect 21821 33269 21833 33303
rect 21867 33300 21879 33303
rect 23658 33300 23664 33312
rect 21867 33272 23664 33300
rect 21867 33269 21879 33272
rect 21821 33263 21879 33269
rect 23658 33260 23664 33272
rect 23716 33260 23722 33312
rect 23753 33303 23811 33309
rect 23753 33269 23765 33303
rect 23799 33300 23811 33303
rect 24394 33300 24400 33312
rect 23799 33272 24400 33300
rect 23799 33269 23811 33272
rect 23753 33263 23811 33269
rect 24394 33260 24400 33272
rect 24452 33260 24458 33312
rect 31294 33260 31300 33312
rect 31352 33300 31358 33312
rect 31573 33303 31631 33309
rect 31573 33300 31585 33303
rect 31352 33272 31585 33300
rect 31352 33260 31358 33272
rect 31573 33269 31585 33272
rect 31619 33269 31631 33303
rect 31726 33300 31754 33340
rect 31846 33328 31852 33380
rect 31904 33368 31910 33380
rect 32784 33368 32812 33399
rect 33870 33396 33876 33408
rect 33928 33396 33934 33448
rect 31904 33340 32812 33368
rect 34333 33371 34391 33377
rect 31904 33328 31910 33340
rect 34333 33337 34345 33371
rect 34379 33368 34391 33371
rect 34790 33368 34796 33380
rect 34379 33340 34796 33368
rect 34379 33337 34391 33340
rect 34333 33331 34391 33337
rect 34790 33328 34796 33340
rect 34848 33328 34854 33380
rect 32582 33300 32588 33312
rect 31726 33272 32588 33300
rect 31573 33263 31631 33269
rect 32582 33260 32588 33272
rect 32640 33260 32646 33312
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 20625 33099 20683 33105
rect 20625 33065 20637 33099
rect 20671 33096 20683 33099
rect 20806 33096 20812 33108
rect 20671 33068 20812 33096
rect 20671 33065 20683 33068
rect 20625 33059 20683 33065
rect 20806 33056 20812 33068
rect 20864 33056 20870 33108
rect 23750 33056 23756 33108
rect 23808 33096 23814 33108
rect 23845 33099 23903 33105
rect 23845 33096 23857 33099
rect 23808 33068 23857 33096
rect 23808 33056 23814 33068
rect 23845 33065 23857 33068
rect 23891 33065 23903 33099
rect 23845 33059 23903 33065
rect 25317 33099 25375 33105
rect 25317 33065 25329 33099
rect 25363 33096 25375 33099
rect 25590 33096 25596 33108
rect 25363 33068 25596 33096
rect 25363 33065 25375 33068
rect 25317 33059 25375 33065
rect 25590 33056 25596 33068
rect 25648 33056 25654 33108
rect 25869 33099 25927 33105
rect 25869 33065 25881 33099
rect 25915 33096 25927 33099
rect 26234 33096 26240 33108
rect 25915 33068 26240 33096
rect 25915 33065 25927 33068
rect 25869 33059 25927 33065
rect 26234 33056 26240 33068
rect 26292 33056 26298 33108
rect 28169 33099 28227 33105
rect 28169 33065 28181 33099
rect 28215 33096 28227 33099
rect 28534 33096 28540 33108
rect 28215 33068 28540 33096
rect 28215 33065 28227 33068
rect 28169 33059 28227 33065
rect 28534 33056 28540 33068
rect 28592 33056 28598 33108
rect 30009 33099 30067 33105
rect 30009 33065 30021 33099
rect 30055 33065 30067 33099
rect 30009 33059 30067 33065
rect 30193 33099 30251 33105
rect 30193 33065 30205 33099
rect 30239 33096 30251 33099
rect 30239 33068 31524 33096
rect 30239 33065 30251 33068
rect 30193 33059 30251 33065
rect 17589 33031 17647 33037
rect 17589 32997 17601 33031
rect 17635 33028 17647 33031
rect 21821 33031 21879 33037
rect 17635 33000 21588 33028
rect 17635 32997 17647 33000
rect 17589 32991 17647 32997
rect 20809 32963 20867 32969
rect 20809 32929 20821 32963
rect 20855 32960 20867 32963
rect 21361 32963 21419 32969
rect 21361 32960 21373 32963
rect 20855 32932 21373 32960
rect 20855 32929 20867 32932
rect 20809 32923 20867 32929
rect 21361 32929 21373 32932
rect 21407 32929 21419 32963
rect 21361 32923 21419 32929
rect 1397 32895 1455 32901
rect 1397 32861 1409 32895
rect 1443 32892 1455 32895
rect 1486 32892 1492 32904
rect 1443 32864 1492 32892
rect 1443 32861 1455 32864
rect 1397 32855 1455 32861
rect 1486 32852 1492 32864
rect 1544 32852 1550 32904
rect 16758 32892 16764 32904
rect 16719 32864 16764 32892
rect 16758 32852 16764 32864
rect 16816 32852 16822 32904
rect 16850 32852 16856 32904
rect 16908 32892 16914 32904
rect 17037 32895 17095 32901
rect 17037 32892 17049 32895
rect 16908 32864 17049 32892
rect 16908 32852 16914 32864
rect 17037 32861 17049 32864
rect 17083 32861 17095 32895
rect 17218 32892 17224 32904
rect 17179 32864 17224 32892
rect 17037 32855 17095 32861
rect 17218 32852 17224 32864
rect 17276 32852 17282 32904
rect 18046 32892 18052 32904
rect 18007 32864 18052 32892
rect 18046 32852 18052 32864
rect 18104 32852 18110 32904
rect 20349 32895 20407 32901
rect 20349 32861 20361 32895
rect 20395 32861 20407 32895
rect 20349 32855 20407 32861
rect 17589 32827 17647 32833
rect 17589 32793 17601 32827
rect 17635 32793 17647 32827
rect 20364 32824 20392 32855
rect 20714 32852 20720 32904
rect 20772 32892 20778 32904
rect 21453 32895 21511 32901
rect 21453 32892 21465 32895
rect 20772 32864 21465 32892
rect 20772 32852 20778 32864
rect 21453 32861 21465 32864
rect 21499 32861 21511 32895
rect 21560 32892 21588 33000
rect 21821 32997 21833 33031
rect 21867 33028 21879 33031
rect 22278 33028 22284 33040
rect 21867 33000 22284 33028
rect 21867 32997 21879 33000
rect 21821 32991 21879 32997
rect 22278 32988 22284 33000
rect 22336 32988 22342 33040
rect 24670 33028 24676 33040
rect 24631 33000 24676 33028
rect 24670 32988 24676 33000
rect 24728 32988 24734 33040
rect 26510 33028 26516 33040
rect 25792 33000 26516 33028
rect 23477 32963 23535 32969
rect 23477 32929 23489 32963
rect 23523 32960 23535 32963
rect 23750 32960 23756 32972
rect 23523 32932 23756 32960
rect 23523 32929 23535 32932
rect 23477 32923 23535 32929
rect 23750 32920 23756 32932
rect 23808 32960 23814 32972
rect 23808 32932 24440 32960
rect 23808 32920 23814 32932
rect 22186 32892 22192 32904
rect 21560 32864 22192 32892
rect 21453 32855 21511 32861
rect 22186 32852 22192 32864
rect 22244 32892 22250 32904
rect 22281 32895 22339 32901
rect 22281 32892 22293 32895
rect 22244 32864 22293 32892
rect 22244 32852 22250 32864
rect 22281 32861 22293 32864
rect 22327 32861 22339 32895
rect 22281 32855 22339 32861
rect 22465 32895 22523 32901
rect 22465 32861 22477 32895
rect 22511 32861 22523 32895
rect 23658 32892 23664 32904
rect 23619 32864 23664 32892
rect 22465 32855 22523 32861
rect 22480 32824 22508 32855
rect 23658 32852 23664 32864
rect 23716 32852 23722 32904
rect 24412 32901 24440 32932
rect 24397 32895 24455 32901
rect 24397 32861 24409 32895
rect 24443 32861 24455 32895
rect 24670 32892 24676 32904
rect 24631 32864 24676 32892
rect 24397 32855 24455 32861
rect 24670 32852 24676 32864
rect 24728 32852 24734 32904
rect 25222 32892 25228 32904
rect 25183 32864 25228 32892
rect 25222 32852 25228 32864
rect 25280 32852 25286 32904
rect 25409 32895 25467 32901
rect 25409 32861 25421 32895
rect 25455 32861 25467 32895
rect 25792 32892 25820 33000
rect 26510 32988 26516 33000
rect 26568 32988 26574 33040
rect 26973 33031 27031 33037
rect 26973 32997 26985 33031
rect 27019 33028 27031 33031
rect 30024 33028 30052 33059
rect 31202 33028 31208 33040
rect 27019 33000 29960 33028
rect 30024 33000 31208 33028
rect 27019 32997 27031 33000
rect 26973 32991 27031 32997
rect 25866 32920 25872 32972
rect 25924 32960 25930 32972
rect 26145 32963 26203 32969
rect 26145 32960 26157 32963
rect 25924 32932 26157 32960
rect 25924 32920 25930 32932
rect 26145 32929 26157 32932
rect 26191 32929 26203 32963
rect 26145 32923 26203 32929
rect 26237 32963 26295 32969
rect 26237 32929 26249 32963
rect 26283 32960 26295 32963
rect 26418 32960 26424 32972
rect 26283 32932 26424 32960
rect 26283 32929 26295 32932
rect 26237 32923 26295 32929
rect 26418 32920 26424 32932
rect 26476 32920 26482 32972
rect 29086 32960 29092 32972
rect 28368 32932 29092 32960
rect 26053 32895 26111 32901
rect 26053 32892 26065 32895
rect 25792 32864 26065 32892
rect 25409 32855 25467 32861
rect 26053 32861 26065 32864
rect 26099 32861 26111 32895
rect 26053 32855 26111 32861
rect 24118 32824 24124 32836
rect 20364 32796 21956 32824
rect 22480 32796 24124 32824
rect 17589 32787 17647 32793
rect 1578 32756 1584 32768
rect 1539 32728 1584 32756
rect 1578 32716 1584 32728
rect 1636 32716 1642 32768
rect 17310 32716 17316 32768
rect 17368 32756 17374 32768
rect 17604 32756 17632 32787
rect 21928 32768 21956 32796
rect 24118 32784 24124 32796
rect 24176 32784 24182 32836
rect 24854 32784 24860 32836
rect 24912 32824 24918 32836
rect 25424 32824 25452 32855
rect 26326 32852 26332 32904
rect 26384 32892 26390 32904
rect 26513 32895 26571 32901
rect 26384 32864 26429 32892
rect 26384 32852 26390 32864
rect 26513 32861 26525 32895
rect 26559 32861 26571 32895
rect 27157 32895 27215 32901
rect 27157 32892 27169 32895
rect 26513 32855 26571 32861
rect 26804 32864 27169 32892
rect 24912 32796 25452 32824
rect 24912 32784 24918 32796
rect 25774 32784 25780 32836
rect 25832 32824 25838 32836
rect 26528 32824 26556 32855
rect 25832 32796 26556 32824
rect 25832 32784 25838 32796
rect 18138 32756 18144 32768
rect 17368 32728 17632 32756
rect 18099 32728 18144 32756
rect 17368 32716 17374 32728
rect 18138 32716 18144 32728
rect 18196 32716 18202 32768
rect 21910 32716 21916 32768
rect 21968 32756 21974 32768
rect 22373 32759 22431 32765
rect 22373 32756 22385 32759
rect 21968 32728 22385 32756
rect 21968 32716 21974 32728
rect 22373 32725 22385 32728
rect 22419 32725 22431 32759
rect 22373 32719 22431 32725
rect 23198 32716 23204 32768
rect 23256 32756 23262 32768
rect 26804 32756 26832 32864
rect 27157 32861 27169 32864
rect 27203 32861 27215 32895
rect 27430 32892 27436 32904
rect 27391 32864 27436 32892
rect 27157 32855 27215 32861
rect 27172 32824 27200 32855
rect 27430 32852 27436 32864
rect 27488 32852 27494 32904
rect 28368 32901 28396 32932
rect 29086 32920 29092 32932
rect 29144 32920 29150 32972
rect 29638 32920 29644 32972
rect 29696 32960 29702 32972
rect 29825 32963 29883 32969
rect 29825 32960 29837 32963
rect 29696 32932 29837 32960
rect 29696 32920 29702 32932
rect 29825 32929 29837 32932
rect 29871 32929 29883 32963
rect 29932 32960 29960 33000
rect 31202 32988 31208 33000
rect 31260 32988 31266 33040
rect 30374 32960 30380 32972
rect 29932 32932 30380 32960
rect 29825 32923 29883 32929
rect 30374 32920 30380 32932
rect 30432 32920 30438 32972
rect 30926 32920 30932 32972
rect 30984 32960 30990 32972
rect 31113 32963 31171 32969
rect 31113 32960 31125 32963
rect 30984 32932 31125 32960
rect 30984 32920 30990 32932
rect 31113 32929 31125 32932
rect 31159 32929 31171 32963
rect 31496 32960 31524 33068
rect 32490 33056 32496 33108
rect 32548 33096 32554 33108
rect 33045 33099 33103 33105
rect 33045 33096 33057 33099
rect 32548 33068 33057 33096
rect 32548 33056 32554 33068
rect 33045 33065 33057 33068
rect 33091 33065 33103 33099
rect 33045 33059 33103 33065
rect 31665 33031 31723 33037
rect 31665 32997 31677 33031
rect 31711 33028 31723 33031
rect 31754 33028 31760 33040
rect 31711 33000 31760 33028
rect 31711 32997 31723 33000
rect 31665 32991 31723 32997
rect 31754 32988 31760 33000
rect 31812 32988 31818 33040
rect 33410 33028 33416 33040
rect 32232 33000 33416 33028
rect 32232 32960 32260 33000
rect 33410 32988 33416 33000
rect 33468 33028 33474 33040
rect 33468 33000 33732 33028
rect 33468 32988 33474 33000
rect 33042 32960 33048 32972
rect 31496 32932 32260 32960
rect 32324 32932 33048 32960
rect 31113 32923 31171 32929
rect 28353 32895 28411 32901
rect 28353 32861 28365 32895
rect 28399 32861 28411 32895
rect 28353 32855 28411 32861
rect 28537 32895 28595 32901
rect 28537 32861 28549 32895
rect 28583 32861 28595 32895
rect 28537 32855 28595 32861
rect 28629 32895 28687 32901
rect 28629 32861 28641 32895
rect 28675 32892 28687 32895
rect 28994 32892 29000 32904
rect 28675 32864 29000 32892
rect 28675 32861 28687 32864
rect 28629 32855 28687 32861
rect 27172 32796 27568 32824
rect 27338 32756 27344 32768
rect 23256 32728 26832 32756
rect 27299 32728 27344 32756
rect 23256 32716 23262 32728
rect 27338 32716 27344 32728
rect 27396 32716 27402 32768
rect 27540 32756 27568 32796
rect 27614 32784 27620 32836
rect 27672 32824 27678 32836
rect 28442 32824 28448 32836
rect 27672 32796 28448 32824
rect 27672 32784 27678 32796
rect 28442 32784 28448 32796
rect 28500 32824 28506 32836
rect 28552 32824 28580 32855
rect 28994 32852 29000 32864
rect 29052 32852 29058 32904
rect 29914 32852 29920 32904
rect 29972 32892 29978 32904
rect 30009 32895 30067 32901
rect 30009 32892 30021 32895
rect 29972 32864 30021 32892
rect 29972 32852 29978 32864
rect 30009 32861 30021 32864
rect 30055 32861 30067 32895
rect 30009 32855 30067 32861
rect 31665 32895 31723 32901
rect 31665 32861 31677 32895
rect 31711 32861 31723 32895
rect 31846 32892 31852 32904
rect 31807 32864 31852 32892
rect 31665 32855 31723 32861
rect 28500 32796 28580 32824
rect 29549 32827 29607 32833
rect 28500 32784 28506 32796
rect 29549 32793 29561 32827
rect 29595 32824 29607 32827
rect 30650 32824 30656 32836
rect 29595 32796 30656 32824
rect 29595 32793 29607 32796
rect 29549 32787 29607 32793
rect 30650 32784 30656 32796
rect 30708 32784 30714 32836
rect 30837 32827 30895 32833
rect 30837 32793 30849 32827
rect 30883 32824 30895 32827
rect 31478 32824 31484 32836
rect 30883 32796 31484 32824
rect 30883 32793 30895 32796
rect 30837 32787 30895 32793
rect 31478 32784 31484 32796
rect 31536 32784 31542 32836
rect 31680 32824 31708 32855
rect 31846 32852 31852 32864
rect 31904 32852 31910 32904
rect 32324 32901 32352 32932
rect 33042 32920 33048 32932
rect 33100 32960 33106 32972
rect 33704 32969 33732 33000
rect 33505 32963 33563 32969
rect 33505 32960 33517 32963
rect 33100 32932 33517 32960
rect 33100 32920 33106 32932
rect 33505 32929 33517 32932
rect 33551 32929 33563 32963
rect 33505 32923 33563 32929
rect 33689 32963 33747 32969
rect 33689 32929 33701 32963
rect 33735 32929 33747 32963
rect 34790 32960 34796 32972
rect 34751 32932 34796 32960
rect 33689 32923 33747 32929
rect 34790 32920 34796 32932
rect 34848 32920 34854 32972
rect 32309 32895 32367 32901
rect 32309 32861 32321 32895
rect 32355 32861 32367 32895
rect 32490 32892 32496 32904
rect 32451 32864 32496 32892
rect 32309 32855 32367 32861
rect 32490 32852 32496 32864
rect 32548 32852 32554 32904
rect 32585 32895 32643 32901
rect 32585 32861 32597 32895
rect 32631 32861 32643 32895
rect 32585 32855 32643 32861
rect 31754 32824 31760 32836
rect 31680 32796 31760 32824
rect 31754 32784 31760 32796
rect 31812 32784 31818 32836
rect 31938 32784 31944 32836
rect 31996 32824 32002 32836
rect 32600 32824 32628 32855
rect 32674 32852 32680 32904
rect 32732 32892 32738 32904
rect 32858 32892 32864 32904
rect 32732 32864 32777 32892
rect 32819 32864 32864 32892
rect 32732 32852 32738 32864
rect 32858 32852 32864 32864
rect 32916 32852 32922 32904
rect 32950 32852 32956 32904
rect 33008 32892 33014 32904
rect 33781 32895 33839 32901
rect 33781 32892 33793 32895
rect 33008 32864 33793 32892
rect 33008 32852 33014 32864
rect 33781 32861 33793 32864
rect 33827 32861 33839 32895
rect 33781 32855 33839 32861
rect 33873 32895 33931 32901
rect 33873 32861 33885 32895
rect 33919 32861 33931 32895
rect 33873 32855 33931 32861
rect 32766 32824 32772 32836
rect 31996 32796 32772 32824
rect 31996 32784 32002 32796
rect 32766 32784 32772 32796
rect 32824 32824 32830 32836
rect 33888 32824 33916 32855
rect 33962 32852 33968 32904
rect 34020 32892 34026 32904
rect 34885 32895 34943 32901
rect 34885 32892 34897 32895
rect 34020 32864 34897 32892
rect 34020 32852 34026 32864
rect 34885 32861 34897 32864
rect 34931 32861 34943 32895
rect 34885 32855 34943 32861
rect 32824 32796 33916 32824
rect 32824 32784 32830 32796
rect 28166 32756 28172 32768
rect 27540 32728 28172 32756
rect 28166 32716 28172 32728
rect 28224 32716 28230 32768
rect 28534 32716 28540 32768
rect 28592 32756 28598 32768
rect 30742 32756 30748 32768
rect 28592 32728 30748 32756
rect 28592 32716 28598 32728
rect 30742 32716 30748 32728
rect 30800 32716 30806 32768
rect 33778 32716 33784 32768
rect 33836 32756 33842 32768
rect 35253 32759 35311 32765
rect 35253 32756 35265 32759
rect 33836 32728 35265 32756
rect 33836 32716 33842 32728
rect 35253 32725 35265 32728
rect 35299 32725 35311 32759
rect 35253 32719 35311 32725
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 16853 32555 16911 32561
rect 16853 32521 16865 32555
rect 16899 32552 16911 32555
rect 18535 32555 18593 32561
rect 16899 32524 18460 32552
rect 16899 32521 16911 32524
rect 16853 32515 16911 32521
rect 18325 32487 18383 32493
rect 17052 32456 17448 32484
rect 15749 32419 15807 32425
rect 15749 32385 15761 32419
rect 15795 32416 15807 32419
rect 16298 32416 16304 32428
rect 15795 32388 16304 32416
rect 15795 32385 15807 32388
rect 15749 32379 15807 32385
rect 16298 32376 16304 32388
rect 16356 32376 16362 32428
rect 16758 32376 16764 32428
rect 16816 32416 16822 32428
rect 17052 32425 17080 32456
rect 17037 32419 17095 32425
rect 17037 32416 17049 32419
rect 16816 32388 17049 32416
rect 16816 32376 16822 32388
rect 17037 32385 17049 32388
rect 17083 32385 17095 32419
rect 17310 32416 17316 32428
rect 17271 32388 17316 32416
rect 17037 32379 17095 32385
rect 17310 32376 17316 32388
rect 17368 32376 17374 32428
rect 15286 32308 15292 32360
rect 15344 32348 15350 32360
rect 15657 32351 15715 32357
rect 15657 32348 15669 32351
rect 15344 32320 15669 32348
rect 15344 32308 15350 32320
rect 15657 32317 15669 32320
rect 15703 32317 15715 32351
rect 17218 32348 17224 32360
rect 15657 32311 15715 32317
rect 16546 32320 17224 32348
rect 16117 32283 16175 32289
rect 16117 32249 16129 32283
rect 16163 32280 16175 32283
rect 16546 32280 16574 32320
rect 17218 32308 17224 32320
rect 17276 32308 17282 32360
rect 17420 32348 17448 32456
rect 18325 32453 18337 32487
rect 18371 32453 18383 32487
rect 18432 32484 18460 32524
rect 18535 32521 18547 32555
rect 18581 32552 18593 32555
rect 19058 32552 19064 32564
rect 18581 32524 19064 32552
rect 18581 32521 18593 32524
rect 18535 32515 18593 32521
rect 19058 32512 19064 32524
rect 19116 32552 19122 32564
rect 19337 32555 19395 32561
rect 19337 32552 19349 32555
rect 19116 32524 19349 32552
rect 19116 32512 19122 32524
rect 19337 32521 19349 32524
rect 19383 32521 19395 32555
rect 19337 32515 19395 32521
rect 21082 32512 21088 32564
rect 21140 32561 21146 32564
rect 21140 32555 21159 32561
rect 21147 32521 21159 32555
rect 21140 32515 21159 32521
rect 23569 32555 23627 32561
rect 23569 32521 23581 32555
rect 23615 32521 23627 32555
rect 23569 32515 23627 32521
rect 21140 32512 21146 32515
rect 20806 32484 20812 32496
rect 18432 32456 20812 32484
rect 18325 32447 18383 32453
rect 17497 32419 17555 32425
rect 17497 32385 17509 32419
rect 17543 32416 17555 32419
rect 18138 32416 18144 32428
rect 17543 32388 18144 32416
rect 17543 32385 17555 32388
rect 17497 32379 17555 32385
rect 18138 32376 18144 32388
rect 18196 32376 18202 32428
rect 18340 32416 18368 32447
rect 20806 32444 20812 32456
rect 20864 32444 20870 32496
rect 20901 32487 20959 32493
rect 20901 32453 20913 32487
rect 20947 32484 20959 32487
rect 22278 32484 22284 32496
rect 20947 32456 22284 32484
rect 20947 32453 20959 32456
rect 20901 32447 20959 32453
rect 22278 32444 22284 32456
rect 22336 32484 22342 32496
rect 23584 32484 23612 32515
rect 23658 32512 23664 32564
rect 23716 32552 23722 32564
rect 24670 32552 24676 32564
rect 23716 32524 24676 32552
rect 23716 32512 23722 32524
rect 24670 32512 24676 32524
rect 24728 32552 24734 32564
rect 25961 32555 26019 32561
rect 24728 32524 25912 32552
rect 24728 32512 24734 32524
rect 22336 32456 23612 32484
rect 24397 32487 24455 32493
rect 22336 32444 22342 32456
rect 24397 32453 24409 32487
rect 24443 32484 24455 32487
rect 25222 32484 25228 32496
rect 24443 32456 25228 32484
rect 24443 32453 24455 32456
rect 24397 32447 24455 32453
rect 18966 32416 18972 32428
rect 18340 32388 18972 32416
rect 18966 32376 18972 32388
rect 19024 32376 19030 32428
rect 19150 32376 19156 32428
rect 19208 32416 19214 32428
rect 19278 32419 19336 32425
rect 19278 32416 19290 32419
rect 19208 32388 19290 32416
rect 19208 32376 19214 32388
rect 19278 32385 19290 32388
rect 19324 32385 19336 32419
rect 22557 32419 22615 32425
rect 22557 32416 22569 32419
rect 19278 32379 19336 32385
rect 21284 32388 22569 32416
rect 19797 32351 19855 32357
rect 19797 32348 19809 32351
rect 17420 32320 19809 32348
rect 19797 32317 19809 32320
rect 19843 32348 19855 32351
rect 19978 32348 19984 32360
rect 19843 32320 19984 32348
rect 19843 32317 19855 32320
rect 19797 32311 19855 32317
rect 19978 32308 19984 32320
rect 20036 32308 20042 32360
rect 16163 32252 16574 32280
rect 16163 32249 16175 32252
rect 16117 32243 16175 32249
rect 16850 32240 16856 32292
rect 16908 32280 16914 32292
rect 17129 32283 17187 32289
rect 17129 32280 17141 32283
rect 16908 32252 17141 32280
rect 16908 32240 16914 32252
rect 17129 32249 17141 32252
rect 17175 32249 17187 32283
rect 19242 32280 19248 32292
rect 17129 32243 17187 32249
rect 18524 32252 19248 32280
rect 18524 32221 18552 32252
rect 19242 32240 19248 32252
rect 19300 32240 19306 32292
rect 21284 32289 21312 32388
rect 22557 32385 22569 32388
rect 22603 32385 22615 32419
rect 22830 32416 22836 32428
rect 22743 32388 22836 32416
rect 22557 32379 22615 32385
rect 22830 32376 22836 32388
rect 22888 32376 22894 32428
rect 23014 32416 23020 32428
rect 22975 32388 23020 32416
rect 23014 32376 23020 32388
rect 23072 32416 23078 32428
rect 23477 32419 23535 32425
rect 23477 32416 23489 32419
rect 23072 32388 23489 32416
rect 23072 32376 23078 32388
rect 23477 32385 23489 32388
rect 23523 32385 23535 32419
rect 23477 32379 23535 32385
rect 23566 32376 23572 32428
rect 23624 32416 23630 32428
rect 25148 32425 25176 32456
rect 25222 32444 25228 32456
rect 25280 32444 25286 32496
rect 23661 32419 23719 32425
rect 23661 32416 23673 32419
rect 23624 32388 23673 32416
rect 23624 32376 23630 32388
rect 23661 32385 23673 32388
rect 23707 32385 23719 32419
rect 23661 32379 23719 32385
rect 24305 32419 24363 32425
rect 24305 32385 24317 32419
rect 24351 32385 24363 32419
rect 24305 32379 24363 32385
rect 24489 32419 24547 32425
rect 24489 32385 24501 32419
rect 24535 32416 24547 32419
rect 25133 32419 25191 32425
rect 24535 32388 25084 32416
rect 24535 32385 24547 32388
rect 24489 32379 24547 32385
rect 22848 32348 22876 32376
rect 23750 32348 23756 32360
rect 22848 32320 23756 32348
rect 23750 32308 23756 32320
rect 23808 32308 23814 32360
rect 21269 32283 21327 32289
rect 21269 32249 21281 32283
rect 21315 32249 21327 32283
rect 21269 32243 21327 32249
rect 22373 32283 22431 32289
rect 22373 32249 22385 32283
rect 22419 32280 22431 32283
rect 24320 32280 24348 32379
rect 24854 32308 24860 32360
rect 24912 32348 24918 32360
rect 24949 32351 25007 32357
rect 24949 32348 24961 32351
rect 24912 32320 24961 32348
rect 24912 32308 24918 32320
rect 24949 32317 24961 32320
rect 24995 32317 25007 32351
rect 25056 32348 25084 32388
rect 25133 32385 25145 32419
rect 25179 32385 25191 32419
rect 25774 32416 25780 32428
rect 25133 32379 25191 32385
rect 25240 32388 25780 32416
rect 25240 32348 25268 32388
rect 25774 32376 25780 32388
rect 25832 32376 25838 32428
rect 25884 32416 25912 32524
rect 25961 32521 25973 32555
rect 26007 32552 26019 32555
rect 26326 32552 26332 32564
rect 26007 32524 26332 32552
rect 26007 32521 26019 32524
rect 25961 32515 26019 32521
rect 26326 32512 26332 32524
rect 26384 32512 26390 32564
rect 27154 32512 27160 32564
rect 27212 32552 27218 32564
rect 28534 32552 28540 32564
rect 27212 32524 28540 32552
rect 27212 32512 27218 32524
rect 28534 32512 28540 32524
rect 28592 32512 28598 32564
rect 28994 32512 29000 32564
rect 29052 32552 29058 32564
rect 29181 32555 29239 32561
rect 29181 32552 29193 32555
rect 29052 32524 29193 32552
rect 29052 32512 29058 32524
rect 29181 32521 29193 32524
rect 29227 32521 29239 32555
rect 31570 32552 31576 32564
rect 29181 32515 29239 32521
rect 30300 32524 31576 32552
rect 27338 32484 27344 32496
rect 26344 32456 27344 32484
rect 26050 32416 26056 32428
rect 25884 32388 26056 32416
rect 26050 32376 26056 32388
rect 26108 32416 26114 32428
rect 26344 32425 26372 32456
rect 27338 32444 27344 32456
rect 27396 32444 27402 32496
rect 30300 32493 30328 32524
rect 31570 32512 31576 32524
rect 31628 32512 31634 32564
rect 31662 32512 31668 32564
rect 31720 32552 31726 32564
rect 31720 32524 32352 32552
rect 31720 32512 31726 32524
rect 30285 32487 30343 32493
rect 30285 32453 30297 32487
rect 30331 32453 30343 32487
rect 30285 32447 30343 32453
rect 30466 32444 30472 32496
rect 30524 32493 30530 32496
rect 30524 32487 30553 32493
rect 30541 32453 30553 32487
rect 30524 32447 30553 32453
rect 30524 32444 30530 32447
rect 31386 32444 31392 32496
rect 31444 32484 31450 32496
rect 31444 32456 32168 32484
rect 31444 32444 31450 32456
rect 26145 32419 26203 32425
rect 26145 32416 26157 32419
rect 26108 32388 26157 32416
rect 26108 32376 26114 32388
rect 26145 32385 26157 32388
rect 26191 32385 26203 32419
rect 26145 32379 26203 32385
rect 26329 32419 26387 32425
rect 26329 32385 26341 32419
rect 26375 32385 26387 32419
rect 26329 32379 26387 32385
rect 26421 32419 26479 32425
rect 26421 32385 26433 32419
rect 26467 32385 26479 32419
rect 26421 32379 26479 32385
rect 25056 32320 25268 32348
rect 24949 32311 25007 32317
rect 25038 32280 25044 32292
rect 22419 32252 25044 32280
rect 22419 32249 22431 32252
rect 22373 32243 22431 32249
rect 25038 32240 25044 32252
rect 25096 32240 25102 32292
rect 26344 32280 26372 32379
rect 25148 32252 26372 32280
rect 26436 32348 26464 32379
rect 26694 32376 26700 32428
rect 26752 32416 26758 32428
rect 27154 32416 27160 32428
rect 26752 32388 27160 32416
rect 26752 32376 26758 32388
rect 27154 32376 27160 32388
rect 27212 32376 27218 32428
rect 27430 32416 27436 32428
rect 27343 32388 27436 32416
rect 27430 32376 27436 32388
rect 27488 32376 27494 32428
rect 28166 32416 28172 32428
rect 28127 32388 28172 32416
rect 28166 32376 28172 32388
rect 28224 32376 28230 32428
rect 28537 32419 28595 32425
rect 28537 32385 28549 32419
rect 28583 32416 28595 32419
rect 29546 32416 29552 32428
rect 28583 32388 29552 32416
rect 28583 32385 28595 32388
rect 28537 32379 28595 32385
rect 29546 32376 29552 32388
rect 29604 32376 29610 32428
rect 30193 32419 30251 32425
rect 30193 32385 30205 32419
rect 30239 32385 30251 32419
rect 30193 32379 30251 32385
rect 27448 32348 27476 32376
rect 26436 32320 27476 32348
rect 18509 32215 18567 32221
rect 18509 32181 18521 32215
rect 18555 32181 18567 32215
rect 18509 32175 18567 32181
rect 18598 32172 18604 32224
rect 18656 32212 18662 32224
rect 18693 32215 18751 32221
rect 18693 32212 18705 32215
rect 18656 32184 18705 32212
rect 18656 32172 18662 32184
rect 18693 32181 18705 32184
rect 18739 32181 18751 32215
rect 18693 32175 18751 32181
rect 19153 32215 19211 32221
rect 19153 32181 19165 32215
rect 19199 32212 19211 32215
rect 19426 32212 19432 32224
rect 19199 32184 19432 32212
rect 19199 32181 19211 32184
rect 19153 32175 19211 32181
rect 19426 32172 19432 32184
rect 19484 32172 19490 32224
rect 19705 32215 19763 32221
rect 19705 32181 19717 32215
rect 19751 32212 19763 32215
rect 20162 32212 20168 32224
rect 19751 32184 20168 32212
rect 19751 32181 19763 32184
rect 19705 32175 19763 32181
rect 20162 32172 20168 32184
rect 20220 32172 20226 32224
rect 21085 32215 21143 32221
rect 21085 32181 21097 32215
rect 21131 32212 21143 32215
rect 21910 32212 21916 32224
rect 21131 32184 21916 32212
rect 21131 32181 21143 32184
rect 21085 32175 21143 32181
rect 21910 32172 21916 32184
rect 21968 32172 21974 32224
rect 24394 32172 24400 32224
rect 24452 32212 24458 32224
rect 25148 32212 25176 32252
rect 25314 32212 25320 32224
rect 24452 32184 25176 32212
rect 25275 32184 25320 32212
rect 24452 32172 24458 32184
rect 25314 32172 25320 32184
rect 25372 32212 25378 32224
rect 26436 32212 26464 32320
rect 28442 32240 28448 32292
rect 28500 32280 28506 32292
rect 30208 32280 30236 32379
rect 30374 32376 30380 32428
rect 30432 32416 30438 32428
rect 31294 32416 31300 32428
rect 30432 32388 30477 32416
rect 31255 32388 31300 32416
rect 30432 32376 30438 32388
rect 31294 32376 31300 32388
rect 31352 32376 31358 32428
rect 31478 32416 31484 32428
rect 31439 32388 31484 32416
rect 31478 32376 31484 32388
rect 31536 32376 31542 32428
rect 32140 32425 32168 32456
rect 32324 32428 32352 32524
rect 32490 32512 32496 32564
rect 32548 32552 32554 32564
rect 33778 32552 33784 32564
rect 32548 32524 32812 32552
rect 33739 32524 33784 32552
rect 32548 32512 32554 32524
rect 32674 32484 32680 32496
rect 32508 32456 32680 32484
rect 32125 32419 32183 32425
rect 32125 32385 32137 32419
rect 32171 32416 32183 32419
rect 32214 32416 32220 32428
rect 32171 32388 32220 32416
rect 32171 32385 32183 32388
rect 32125 32379 32183 32385
rect 32214 32376 32220 32388
rect 32272 32376 32278 32428
rect 32306 32376 32312 32428
rect 32364 32416 32370 32428
rect 32364 32388 32457 32416
rect 32364 32376 32370 32388
rect 30558 32308 30564 32360
rect 30616 32348 30622 32360
rect 30653 32351 30711 32357
rect 30653 32348 30665 32351
rect 30616 32320 30665 32348
rect 30616 32308 30622 32320
rect 30653 32317 30665 32320
rect 30699 32317 30711 32351
rect 30653 32311 30711 32317
rect 30926 32308 30932 32360
rect 30984 32348 30990 32360
rect 30984 32320 31248 32348
rect 30984 32308 30990 32320
rect 31018 32280 31024 32292
rect 28500 32252 30144 32280
rect 30208 32252 31024 32280
rect 28500 32240 28506 32252
rect 26970 32212 26976 32224
rect 25372 32184 26464 32212
rect 26931 32184 26976 32212
rect 25372 32172 25378 32184
rect 26970 32172 26976 32184
rect 27028 32172 27034 32224
rect 28902 32172 28908 32224
rect 28960 32212 28966 32224
rect 30009 32215 30067 32221
rect 30009 32212 30021 32215
rect 28960 32184 30021 32212
rect 28960 32172 28966 32184
rect 30009 32181 30021 32184
rect 30055 32181 30067 32215
rect 30116 32212 30144 32252
rect 31018 32240 31024 32252
rect 31076 32240 31082 32292
rect 30190 32212 30196 32224
rect 30116 32184 30196 32212
rect 30009 32175 30067 32181
rect 30190 32172 30196 32184
rect 30248 32172 30254 32224
rect 31110 32212 31116 32224
rect 31071 32184 31116 32212
rect 31110 32172 31116 32184
rect 31168 32172 31174 32224
rect 31220 32212 31248 32320
rect 31570 32308 31576 32360
rect 31628 32348 31634 32360
rect 31754 32348 31760 32360
rect 31628 32320 31760 32348
rect 31628 32308 31634 32320
rect 31754 32308 31760 32320
rect 31812 32348 31818 32360
rect 32508 32348 32536 32456
rect 32674 32444 32680 32456
rect 32732 32444 32738 32496
rect 32784 32484 32812 32524
rect 33778 32512 33784 32524
rect 33836 32512 33842 32564
rect 33502 32484 33508 32496
rect 32784 32456 33508 32484
rect 33502 32444 33508 32456
rect 33560 32484 33566 32496
rect 33689 32487 33747 32493
rect 33689 32484 33701 32487
rect 33560 32456 33701 32484
rect 33560 32444 33566 32456
rect 33689 32453 33701 32456
rect 33735 32484 33747 32487
rect 33870 32484 33876 32496
rect 33735 32456 33876 32484
rect 33735 32453 33747 32456
rect 33689 32447 33747 32453
rect 33870 32444 33876 32456
rect 33928 32444 33934 32496
rect 32585 32419 32643 32425
rect 32585 32385 32597 32419
rect 32631 32416 32643 32419
rect 32631 32388 33916 32416
rect 32631 32385 32643 32388
rect 32585 32379 32643 32385
rect 31812 32320 32536 32348
rect 31812 32308 31818 32320
rect 31478 32240 31484 32292
rect 31536 32280 31542 32292
rect 32600 32280 32628 32379
rect 33888 32357 33916 32388
rect 32677 32351 32735 32357
rect 32677 32317 32689 32351
rect 32723 32317 32735 32351
rect 32677 32311 32735 32317
rect 33873 32351 33931 32357
rect 33873 32317 33885 32351
rect 33919 32317 33931 32351
rect 33873 32311 33931 32317
rect 31536 32252 32628 32280
rect 32692 32280 32720 32311
rect 34698 32280 34704 32292
rect 32692 32252 34704 32280
rect 31536 32240 31542 32252
rect 34698 32240 34704 32252
rect 34756 32240 34762 32292
rect 31754 32212 31760 32224
rect 31220 32184 31760 32212
rect 31754 32172 31760 32184
rect 31812 32172 31818 32224
rect 33318 32212 33324 32224
rect 33279 32184 33324 32212
rect 33318 32172 33324 32184
rect 33376 32172 33382 32224
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 15286 32008 15292 32020
rect 15247 31980 15292 32008
rect 15286 31968 15292 31980
rect 15344 31968 15350 32020
rect 16298 32008 16304 32020
rect 16259 31980 16304 32008
rect 16298 31968 16304 31980
rect 16356 31968 16362 32020
rect 16945 32011 17003 32017
rect 16945 31977 16957 32011
rect 16991 32008 17003 32011
rect 17310 32008 17316 32020
rect 16991 31980 17316 32008
rect 16991 31977 17003 31980
rect 16945 31971 17003 31977
rect 17310 31968 17316 31980
rect 17368 31968 17374 32020
rect 20346 31968 20352 32020
rect 20404 32008 20410 32020
rect 20625 32011 20683 32017
rect 20625 32008 20637 32011
rect 20404 31980 20637 32008
rect 20404 31968 20410 31980
rect 20625 31977 20637 31980
rect 20671 31977 20683 32011
rect 23198 32008 23204 32020
rect 23159 31980 23204 32008
rect 20625 31971 20683 31977
rect 23198 31968 23204 31980
rect 23256 31968 23262 32020
rect 24765 32011 24823 32017
rect 24765 31977 24777 32011
rect 24811 32008 24823 32011
rect 25314 32008 25320 32020
rect 24811 31980 25320 32008
rect 24811 31977 24823 31980
rect 24765 31971 24823 31977
rect 25314 31968 25320 31980
rect 25372 31968 25378 32020
rect 25682 31968 25688 32020
rect 25740 32008 25746 32020
rect 26510 32008 26516 32020
rect 25740 31980 26516 32008
rect 25740 31968 25746 31980
rect 26510 31968 26516 31980
rect 26568 32008 26574 32020
rect 26881 32011 26939 32017
rect 26881 32008 26893 32011
rect 26568 31980 26893 32008
rect 26568 31968 26574 31980
rect 26881 31977 26893 31980
rect 26927 31977 26939 32011
rect 26881 31971 26939 31977
rect 26970 31968 26976 32020
rect 27028 32008 27034 32020
rect 32950 32008 32956 32020
rect 27028 31980 32956 32008
rect 27028 31968 27034 31980
rect 32950 31968 32956 31980
rect 33008 31968 33014 32020
rect 33502 32008 33508 32020
rect 33463 31980 33508 32008
rect 33502 31968 33508 31980
rect 33560 31968 33566 32020
rect 35618 32008 35624 32020
rect 33612 31980 35624 32008
rect 18509 31943 18567 31949
rect 18509 31940 18521 31943
rect 15948 31912 18521 31940
rect 15654 31832 15660 31884
rect 15712 31872 15718 31884
rect 15948 31881 15976 31912
rect 18509 31909 18521 31912
rect 18555 31940 18567 31943
rect 18782 31940 18788 31952
rect 18555 31912 18788 31940
rect 18555 31909 18567 31912
rect 18509 31903 18567 31909
rect 18782 31900 18788 31912
rect 18840 31900 18846 31952
rect 21082 31900 21088 31952
rect 21140 31940 21146 31952
rect 24949 31943 25007 31949
rect 21140 31912 21772 31940
rect 21140 31900 21146 31912
rect 15933 31875 15991 31881
rect 15933 31872 15945 31875
rect 15712 31844 15945 31872
rect 15712 31832 15718 31844
rect 15933 31841 15945 31844
rect 15979 31841 15991 31875
rect 15933 31835 15991 31841
rect 16206 31832 16212 31884
rect 16264 31872 16270 31884
rect 17037 31875 17095 31881
rect 17037 31872 17049 31875
rect 16264 31844 17049 31872
rect 16264 31832 16270 31844
rect 17037 31841 17049 31844
rect 17083 31841 17095 31875
rect 17037 31835 17095 31841
rect 18233 31875 18291 31881
rect 18233 31841 18245 31875
rect 18279 31872 18291 31875
rect 18598 31872 18604 31884
rect 18279 31844 18604 31872
rect 18279 31841 18291 31844
rect 18233 31835 18291 31841
rect 18598 31832 18604 31844
rect 18656 31832 18662 31884
rect 21744 31881 21772 31912
rect 24949 31909 24961 31943
rect 24995 31940 25007 31943
rect 25038 31940 25044 31952
rect 24995 31912 25044 31940
rect 24995 31909 25007 31912
rect 24949 31903 25007 31909
rect 25038 31900 25044 31912
rect 25096 31900 25102 31952
rect 25593 31943 25651 31949
rect 25593 31909 25605 31943
rect 25639 31940 25651 31943
rect 28629 31943 28687 31949
rect 25639 31912 28580 31940
rect 25639 31909 25651 31912
rect 25593 31903 25651 31909
rect 18693 31875 18751 31881
rect 18693 31841 18705 31875
rect 18739 31872 18751 31875
rect 19337 31875 19395 31881
rect 19337 31872 19349 31875
rect 18739 31844 19349 31872
rect 18739 31841 18751 31844
rect 18693 31835 18751 31841
rect 19337 31841 19349 31844
rect 19383 31841 19395 31875
rect 19337 31835 19395 31841
rect 21729 31875 21787 31881
rect 21729 31841 21741 31875
rect 21775 31841 21787 31875
rect 22278 31872 22284 31884
rect 22239 31844 22284 31872
rect 21729 31835 21787 31841
rect 22278 31832 22284 31844
rect 22336 31832 22342 31884
rect 23661 31875 23719 31881
rect 23661 31841 23673 31875
rect 23707 31872 23719 31875
rect 24578 31872 24584 31884
rect 23707 31844 24584 31872
rect 23707 31841 23719 31844
rect 23661 31835 23719 31841
rect 24578 31832 24584 31844
rect 24636 31832 24642 31884
rect 26053 31875 26111 31881
rect 26053 31841 26065 31875
rect 26099 31872 26111 31875
rect 27522 31872 27528 31884
rect 26099 31844 27528 31872
rect 26099 31841 26111 31844
rect 26053 31835 26111 31841
rect 27522 31832 27528 31844
rect 27580 31832 27586 31884
rect 15289 31807 15347 31813
rect 15289 31773 15301 31807
rect 15335 31773 15347 31807
rect 15470 31804 15476 31816
rect 15431 31776 15476 31804
rect 15289 31767 15347 31773
rect 15304 31736 15332 31767
rect 15470 31764 15476 31776
rect 15528 31764 15534 31816
rect 16117 31807 16175 31813
rect 16117 31773 16129 31807
rect 16163 31773 16175 31807
rect 16758 31804 16764 31816
rect 16719 31776 16764 31804
rect 16117 31767 16175 31773
rect 16022 31736 16028 31748
rect 15304 31708 16028 31736
rect 16022 31696 16028 31708
rect 16080 31696 16086 31748
rect 15930 31628 15936 31680
rect 15988 31668 15994 31680
rect 16132 31668 16160 31767
rect 16758 31764 16764 31776
rect 16816 31764 16822 31816
rect 16850 31764 16856 31816
rect 16908 31804 16914 31816
rect 19426 31804 19432 31816
rect 16908 31776 17724 31804
rect 19387 31776 19432 31804
rect 16908 31764 16914 31776
rect 17034 31696 17040 31748
rect 17092 31736 17098 31748
rect 17589 31739 17647 31745
rect 17589 31736 17601 31739
rect 17092 31708 17601 31736
rect 17092 31696 17098 31708
rect 17589 31705 17601 31708
rect 17635 31705 17647 31739
rect 17696 31736 17724 31776
rect 19426 31764 19432 31776
rect 19484 31764 19490 31816
rect 20809 31807 20867 31813
rect 20809 31773 20821 31807
rect 20855 31773 20867 31807
rect 21082 31804 21088 31816
rect 21043 31776 21088 31804
rect 20809 31767 20867 31773
rect 20162 31736 20168 31748
rect 17696 31708 20168 31736
rect 17589 31699 17647 31705
rect 20162 31696 20168 31708
rect 20220 31696 20226 31748
rect 20824 31736 20852 31767
rect 21082 31764 21088 31776
rect 21140 31764 21146 31816
rect 21910 31804 21916 31816
rect 21871 31776 21916 31804
rect 21910 31764 21916 31776
rect 21968 31764 21974 31816
rect 26142 31804 26148 31816
rect 26103 31776 26148 31804
rect 26142 31764 26148 31776
rect 26200 31764 26206 31816
rect 26789 31807 26847 31813
rect 26789 31804 26801 31807
rect 26252 31776 26801 31804
rect 23750 31736 23756 31748
rect 20824 31708 21956 31736
rect 23711 31708 23756 31736
rect 21928 31680 21956 31708
rect 23750 31696 23756 31708
rect 23808 31696 23814 31748
rect 24394 31696 24400 31748
rect 24452 31736 24458 31748
rect 24581 31739 24639 31745
rect 24581 31736 24593 31739
rect 24452 31708 24593 31736
rect 24452 31696 24458 31708
rect 24581 31705 24593 31708
rect 24627 31705 24639 31739
rect 24581 31699 24639 31705
rect 25958 31696 25964 31748
rect 26016 31736 26022 31748
rect 26252 31736 26280 31776
rect 26789 31773 26801 31776
rect 26835 31773 26847 31807
rect 26789 31767 26847 31773
rect 28166 31764 28172 31816
rect 28224 31804 28230 31816
rect 28261 31807 28319 31813
rect 28261 31804 28273 31807
rect 28224 31776 28273 31804
rect 28224 31764 28230 31776
rect 28261 31773 28273 31776
rect 28307 31773 28319 31807
rect 28442 31804 28448 31816
rect 28403 31776 28448 31804
rect 28261 31767 28319 31773
rect 28442 31764 28448 31776
rect 28500 31764 28506 31816
rect 28552 31804 28580 31912
rect 28629 31909 28641 31943
rect 28675 31940 28687 31943
rect 29086 31940 29092 31952
rect 28675 31912 29092 31940
rect 28675 31909 28687 31912
rect 28629 31903 28687 31909
rect 29086 31900 29092 31912
rect 29144 31900 29150 31952
rect 31570 31940 31576 31952
rect 29472 31912 31576 31940
rect 29472 31804 29500 31912
rect 29546 31832 29552 31884
rect 29604 31872 29610 31884
rect 30558 31872 30564 31884
rect 29604 31844 29649 31872
rect 29748 31844 30564 31872
rect 29604 31832 29610 31844
rect 29748 31804 29776 31844
rect 30558 31832 30564 31844
rect 30616 31832 30622 31884
rect 28552 31776 29500 31804
rect 29656 31776 29776 31804
rect 29825 31807 29883 31813
rect 26016 31708 26280 31736
rect 27617 31739 27675 31745
rect 26016 31696 26022 31708
rect 27617 31705 27629 31739
rect 27663 31705 27675 31739
rect 27617 31699 27675 31705
rect 27801 31739 27859 31745
rect 27801 31705 27813 31739
rect 27847 31736 27859 31739
rect 28534 31736 28540 31748
rect 27847 31708 28540 31736
rect 27847 31705 27859 31708
rect 27801 31699 27859 31705
rect 15988 31640 16160 31668
rect 17681 31671 17739 31677
rect 15988 31628 15994 31640
rect 17681 31637 17693 31671
rect 17727 31668 17739 31671
rect 18046 31668 18052 31680
rect 17727 31640 18052 31668
rect 17727 31637 17739 31640
rect 17681 31631 17739 31637
rect 18046 31628 18052 31640
rect 18104 31668 18110 31680
rect 18230 31668 18236 31680
rect 18104 31640 18236 31668
rect 18104 31628 18110 31640
rect 18230 31628 18236 31640
rect 18288 31628 18294 31680
rect 19426 31628 19432 31680
rect 19484 31668 19490 31680
rect 19797 31671 19855 31677
rect 19797 31668 19809 31671
rect 19484 31640 19809 31668
rect 19484 31628 19490 31640
rect 19797 31637 19809 31640
rect 19843 31637 19855 31671
rect 19797 31631 19855 31637
rect 20714 31628 20720 31680
rect 20772 31668 20778 31680
rect 20993 31671 21051 31677
rect 20993 31668 21005 31671
rect 20772 31640 21005 31668
rect 20772 31628 20778 31640
rect 20993 31637 21005 31640
rect 21039 31668 21051 31671
rect 21818 31668 21824 31680
rect 21039 31640 21824 31668
rect 21039 31637 21051 31640
rect 20993 31631 21051 31637
rect 21818 31628 21824 31640
rect 21876 31628 21882 31680
rect 21910 31628 21916 31680
rect 21968 31628 21974 31680
rect 22189 31671 22247 31677
rect 22189 31637 22201 31671
rect 22235 31668 22247 31671
rect 23382 31668 23388 31680
rect 22235 31640 23388 31668
rect 22235 31637 22247 31640
rect 22189 31631 22247 31637
rect 23382 31628 23388 31640
rect 23440 31628 23446 31680
rect 23474 31628 23480 31680
rect 23532 31668 23538 31680
rect 23661 31671 23719 31677
rect 23661 31668 23673 31671
rect 23532 31640 23673 31668
rect 23532 31628 23538 31640
rect 23661 31637 23673 31640
rect 23707 31637 23719 31671
rect 23661 31631 23719 31637
rect 23842 31628 23848 31680
rect 23900 31668 23906 31680
rect 24781 31671 24839 31677
rect 24781 31668 24793 31671
rect 23900 31640 24793 31668
rect 23900 31628 23906 31640
rect 24781 31637 24793 31640
rect 24827 31637 24839 31671
rect 24781 31631 24839 31637
rect 25682 31628 25688 31680
rect 25740 31668 25746 31680
rect 26053 31671 26111 31677
rect 26053 31668 26065 31671
rect 25740 31640 26065 31668
rect 25740 31628 25746 31640
rect 26053 31637 26065 31640
rect 26099 31637 26111 31671
rect 27632 31668 27660 31699
rect 28534 31696 28540 31708
rect 28592 31736 28598 31748
rect 29656 31736 29684 31776
rect 29825 31773 29837 31807
rect 29871 31804 29883 31807
rect 30190 31804 30196 31816
rect 29871 31776 30196 31804
rect 29871 31773 29883 31776
rect 29825 31767 29883 31773
rect 30190 31764 30196 31776
rect 30248 31764 30254 31816
rect 30668 31804 30696 31912
rect 31570 31900 31576 31912
rect 31628 31900 31634 31952
rect 32582 31900 32588 31952
rect 32640 31940 32646 31952
rect 33612 31940 33640 31980
rect 35618 31968 35624 31980
rect 35676 31968 35682 32020
rect 34146 31940 34152 31952
rect 32640 31912 33640 31940
rect 33704 31912 34152 31940
rect 32640 31900 32646 31912
rect 30926 31832 30932 31884
rect 30984 31872 30990 31884
rect 33042 31872 33048 31884
rect 30984 31844 31340 31872
rect 30984 31832 30990 31844
rect 31312 31813 31340 31844
rect 32508 31844 33048 31872
rect 31205 31807 31263 31813
rect 31205 31804 31217 31807
rect 30668 31776 31217 31804
rect 31205 31773 31217 31776
rect 31251 31773 31263 31807
rect 31205 31767 31263 31773
rect 31297 31807 31355 31813
rect 31297 31773 31309 31807
rect 31343 31773 31355 31807
rect 31297 31767 31355 31773
rect 31386 31764 31392 31816
rect 31444 31804 31450 31816
rect 31573 31807 31631 31813
rect 31444 31776 31489 31804
rect 31444 31764 31450 31776
rect 31573 31773 31585 31807
rect 31619 31773 31631 31807
rect 32214 31804 32220 31816
rect 32175 31776 32220 31804
rect 31573 31767 31631 31773
rect 28592 31708 29684 31736
rect 28592 31696 28598 31708
rect 31478 31696 31484 31748
rect 31536 31736 31542 31748
rect 31588 31736 31616 31767
rect 32214 31764 32220 31776
rect 32272 31764 32278 31816
rect 32306 31764 32312 31816
rect 32364 31804 32370 31816
rect 32508 31813 32536 31844
rect 33042 31832 33048 31844
rect 33100 31832 33106 31884
rect 33226 31832 33232 31884
rect 33284 31872 33290 31884
rect 33704 31872 33732 31912
rect 34146 31900 34152 31912
rect 34204 31900 34210 31952
rect 34698 31900 34704 31952
rect 34756 31940 34762 31952
rect 36078 31940 36084 31952
rect 34756 31912 36084 31940
rect 34756 31900 34762 31912
rect 36078 31900 36084 31912
rect 36136 31900 36142 31952
rect 33284 31844 33732 31872
rect 34057 31875 34115 31881
rect 33284 31832 33290 31844
rect 34057 31841 34069 31875
rect 34103 31872 34115 31875
rect 35526 31872 35532 31884
rect 34103 31844 35532 31872
rect 34103 31841 34115 31844
rect 34057 31835 34115 31841
rect 35526 31832 35532 31844
rect 35584 31832 35590 31884
rect 32493 31807 32551 31813
rect 32364 31776 32409 31804
rect 32364 31764 32370 31776
rect 32493 31773 32505 31807
rect 32539 31773 32551 31807
rect 32493 31767 32551 31773
rect 32582 31764 32588 31816
rect 32640 31804 32646 31816
rect 32640 31776 32685 31804
rect 32640 31764 32646 31776
rect 32950 31764 32956 31816
rect 33008 31804 33014 31816
rect 33137 31807 33195 31813
rect 33137 31804 33149 31807
rect 33008 31776 33149 31804
rect 33008 31764 33014 31776
rect 33137 31773 33149 31776
rect 33183 31773 33195 31807
rect 33137 31767 33195 31773
rect 33321 31807 33379 31813
rect 33321 31773 33333 31807
rect 33367 31804 33379 31807
rect 33410 31804 33416 31816
rect 33367 31776 33416 31804
rect 33367 31773 33379 31776
rect 33321 31767 33379 31773
rect 33410 31764 33416 31776
rect 33468 31764 33474 31816
rect 33965 31807 34023 31813
rect 33520 31801 33916 31804
rect 33965 31801 33977 31807
rect 33520 31776 33977 31801
rect 31536 31708 31616 31736
rect 31536 31696 31542 31708
rect 31846 31696 31852 31748
rect 31904 31736 31910 31748
rect 33520 31736 33548 31776
rect 33888 31773 33977 31776
rect 34011 31773 34023 31807
rect 34146 31804 34152 31816
rect 34107 31776 34152 31804
rect 33965 31767 34023 31773
rect 34146 31764 34152 31776
rect 34204 31764 34210 31816
rect 34698 31804 34704 31816
rect 34659 31776 34704 31804
rect 34698 31764 34704 31776
rect 34756 31764 34762 31816
rect 34885 31807 34943 31813
rect 34885 31804 34897 31807
rect 34808 31776 34897 31804
rect 31904 31708 33548 31736
rect 31904 31696 31910 31708
rect 34054 31696 34060 31748
rect 34112 31736 34118 31748
rect 34808 31736 34836 31776
rect 34885 31773 34897 31776
rect 34931 31773 34943 31807
rect 34885 31767 34943 31773
rect 34112 31708 34836 31736
rect 34112 31696 34118 31708
rect 28718 31668 28724 31680
rect 27632 31640 28724 31668
rect 26053 31631 26111 31637
rect 28718 31628 28724 31640
rect 28776 31628 28782 31680
rect 30929 31671 30987 31677
rect 30929 31637 30941 31671
rect 30975 31668 30987 31671
rect 31570 31668 31576 31680
rect 30975 31640 31576 31668
rect 30975 31637 30987 31640
rect 30929 31631 30987 31637
rect 31570 31628 31576 31640
rect 31628 31628 31634 31680
rect 32030 31668 32036 31680
rect 31991 31640 32036 31668
rect 32030 31628 32036 31640
rect 32088 31628 32094 31680
rect 34514 31628 34520 31680
rect 34572 31668 34578 31680
rect 34793 31671 34851 31677
rect 34793 31668 34805 31671
rect 34572 31640 34805 31668
rect 34572 31628 34578 31640
rect 34793 31637 34805 31640
rect 34839 31637 34851 31671
rect 34793 31631 34851 31637
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 15197 31467 15255 31473
rect 15197 31433 15209 31467
rect 15243 31464 15255 31467
rect 15470 31464 15476 31476
rect 15243 31436 15476 31464
rect 15243 31433 15255 31436
rect 15197 31427 15255 31433
rect 15470 31424 15476 31436
rect 15528 31424 15534 31476
rect 16022 31424 16028 31476
rect 16080 31464 16086 31476
rect 16117 31467 16175 31473
rect 16117 31464 16129 31467
rect 16080 31436 16129 31464
rect 16080 31424 16086 31436
rect 16117 31433 16129 31436
rect 16163 31433 16175 31467
rect 16850 31464 16856 31476
rect 16811 31436 16856 31464
rect 16117 31427 16175 31433
rect 16132 31396 16160 31427
rect 16850 31424 16856 31436
rect 16908 31424 16914 31476
rect 18322 31464 18328 31476
rect 18283 31436 18328 31464
rect 18322 31424 18328 31436
rect 18380 31424 18386 31476
rect 18782 31464 18788 31476
rect 18743 31436 18788 31464
rect 18782 31424 18788 31436
rect 18840 31424 18846 31476
rect 19153 31467 19211 31473
rect 19153 31433 19165 31467
rect 19199 31464 19211 31467
rect 19242 31464 19248 31476
rect 19199 31436 19248 31464
rect 19199 31433 19211 31436
rect 19153 31427 19211 31433
rect 19242 31424 19248 31436
rect 19300 31424 19306 31476
rect 19334 31424 19340 31476
rect 19392 31464 19398 31476
rect 19392 31436 20199 31464
rect 19392 31424 19398 31436
rect 17957 31399 18015 31405
rect 15120 31368 15976 31396
rect 16132 31368 17172 31396
rect 15120 31337 15148 31368
rect 15105 31331 15163 31337
rect 15105 31297 15117 31331
rect 15151 31297 15163 31331
rect 15286 31328 15292 31340
rect 15247 31300 15292 31328
rect 15105 31291 15163 31297
rect 15286 31288 15292 31300
rect 15344 31288 15350 31340
rect 15948 31337 15976 31368
rect 15933 31331 15991 31337
rect 15933 31297 15945 31331
rect 15979 31328 15991 31331
rect 16022 31328 16028 31340
rect 15979 31300 16028 31328
rect 15979 31297 15991 31300
rect 15933 31291 15991 31297
rect 16022 31288 16028 31300
rect 16080 31288 16086 31340
rect 16850 31288 16856 31340
rect 16908 31328 16914 31340
rect 17034 31328 17040 31340
rect 16908 31300 17040 31328
rect 16908 31288 16914 31300
rect 17034 31288 17040 31300
rect 17092 31288 17098 31340
rect 17144 31337 17172 31368
rect 17957 31365 17969 31399
rect 18003 31365 18015 31399
rect 17957 31359 18015 31365
rect 18173 31399 18231 31405
rect 18173 31365 18185 31399
rect 18219 31396 18231 31399
rect 19426 31396 19432 31408
rect 18219 31368 19432 31396
rect 18219 31365 18231 31368
rect 18173 31359 18231 31365
rect 17129 31331 17187 31337
rect 17129 31297 17141 31331
rect 17175 31297 17187 31331
rect 17129 31291 17187 31297
rect 17313 31331 17371 31337
rect 17313 31297 17325 31331
rect 17359 31328 17371 31331
rect 17862 31328 17868 31340
rect 17359 31300 17868 31328
rect 17359 31297 17371 31300
rect 17313 31291 17371 31297
rect 15749 31263 15807 31269
rect 15749 31229 15761 31263
rect 15795 31260 15807 31263
rect 15838 31260 15844 31272
rect 15795 31232 15844 31260
rect 15795 31229 15807 31232
rect 15749 31223 15807 31229
rect 15838 31220 15844 31232
rect 15896 31220 15902 31272
rect 17144 31260 17172 31291
rect 17862 31288 17868 31300
rect 17920 31288 17926 31340
rect 17972 31328 18000 31359
rect 19426 31356 19432 31368
rect 19484 31356 19490 31408
rect 20171 31396 20199 31436
rect 20254 31424 20260 31476
rect 20312 31464 20318 31476
rect 21821 31467 21879 31473
rect 21821 31464 21833 31467
rect 20312 31436 21833 31464
rect 20312 31424 20318 31436
rect 21821 31433 21833 31436
rect 21867 31433 21879 31467
rect 24578 31464 24584 31476
rect 24539 31436 24584 31464
rect 21821 31427 21879 31433
rect 24578 31424 24584 31436
rect 24636 31424 24642 31476
rect 26786 31424 26792 31476
rect 26844 31464 26850 31476
rect 26844 31436 27108 31464
rect 26844 31424 26850 31436
rect 21085 31399 21143 31405
rect 21085 31396 21097 31399
rect 20171 31368 21097 31396
rect 18506 31328 18512 31340
rect 17972 31300 18512 31328
rect 18506 31288 18512 31300
rect 18564 31288 18570 31340
rect 18966 31328 18972 31340
rect 18879 31300 18972 31328
rect 18966 31288 18972 31300
rect 19024 31328 19030 31340
rect 19024 31300 19104 31328
rect 19024 31288 19030 31300
rect 17954 31260 17960 31272
rect 17144 31232 17960 31260
rect 17954 31220 17960 31232
rect 18012 31220 18018 31272
rect 15194 31152 15200 31204
rect 15252 31192 15258 31204
rect 17221 31195 17279 31201
rect 17221 31192 17233 31195
rect 15252 31164 17233 31192
rect 15252 31152 15258 31164
rect 17221 31161 17233 31164
rect 17267 31192 17279 31195
rect 18046 31192 18052 31204
rect 17267 31164 18052 31192
rect 17267 31161 17279 31164
rect 17221 31155 17279 31161
rect 18046 31152 18052 31164
rect 18104 31152 18110 31204
rect 19076 31192 19104 31300
rect 19150 31288 19156 31340
rect 19208 31328 19214 31340
rect 19245 31331 19303 31337
rect 19245 31328 19257 31331
rect 19208 31300 19257 31328
rect 19208 31288 19214 31300
rect 19245 31297 19257 31300
rect 19291 31297 19303 31331
rect 20070 31328 20076 31340
rect 20031 31300 20076 31328
rect 19245 31291 19303 31297
rect 20070 31288 20076 31300
rect 20128 31288 20134 31340
rect 20171 31328 20199 31368
rect 21085 31365 21097 31368
rect 21131 31365 21143 31399
rect 24670 31396 24676 31408
rect 21085 31359 21143 31365
rect 23860 31368 24676 31396
rect 20349 31331 20407 31337
rect 20349 31328 20361 31331
rect 20171 31300 20361 31328
rect 20349 31297 20361 31300
rect 20395 31297 20407 31331
rect 20349 31291 20407 31297
rect 20993 31331 21051 31337
rect 20993 31297 21005 31331
rect 21039 31297 21051 31331
rect 21174 31328 21180 31340
rect 21135 31300 21180 31328
rect 20993 31291 21051 31297
rect 20162 31260 20168 31272
rect 20123 31232 20168 31260
rect 20162 31220 20168 31232
rect 20220 31220 20226 31272
rect 20254 31192 20260 31204
rect 19076 31164 20260 31192
rect 20254 31152 20260 31164
rect 20312 31152 20318 31204
rect 20533 31195 20591 31201
rect 20533 31161 20545 31195
rect 20579 31192 20591 31195
rect 20714 31192 20720 31204
rect 20579 31164 20720 31192
rect 20579 31161 20591 31164
rect 20533 31155 20591 31161
rect 20714 31152 20720 31164
rect 20772 31152 20778 31204
rect 21008 31192 21036 31291
rect 21174 31288 21180 31300
rect 21232 31288 21238 31340
rect 21818 31288 21824 31340
rect 21876 31328 21882 31340
rect 22097 31331 22155 31337
rect 22097 31328 22109 31331
rect 21876 31300 22109 31328
rect 21876 31288 21882 31300
rect 22097 31297 22109 31300
rect 22143 31297 22155 31331
rect 22097 31291 22155 31297
rect 23017 31331 23075 31337
rect 23017 31297 23029 31331
rect 23063 31328 23075 31331
rect 23106 31328 23112 31340
rect 23063 31300 23112 31328
rect 23063 31297 23075 31300
rect 23017 31291 23075 31297
rect 23106 31288 23112 31300
rect 23164 31288 23170 31340
rect 23860 31337 23888 31368
rect 24670 31356 24676 31368
rect 24728 31356 24734 31408
rect 26050 31356 26056 31408
rect 26108 31396 26114 31408
rect 26108 31368 27016 31396
rect 26108 31356 26114 31368
rect 23845 31331 23903 31337
rect 23845 31297 23857 31331
rect 23891 31297 23903 31331
rect 24026 31328 24032 31340
rect 23987 31300 24032 31328
rect 23845 31291 23903 31297
rect 24026 31288 24032 31300
rect 24084 31288 24090 31340
rect 24489 31331 24547 31337
rect 24489 31297 24501 31331
rect 24535 31297 24547 31331
rect 24489 31291 24547 31297
rect 21082 31220 21088 31272
rect 21140 31260 21146 31272
rect 22002 31260 22008 31272
rect 21140 31232 22008 31260
rect 21140 31220 21146 31232
rect 22002 31220 22008 31232
rect 22060 31220 22066 31272
rect 22189 31263 22247 31269
rect 22189 31229 22201 31263
rect 22235 31229 22247 31263
rect 22189 31223 22247 31229
rect 22281 31263 22339 31269
rect 22281 31229 22293 31263
rect 22327 31229 22339 31263
rect 22281 31223 22339 31229
rect 21450 31192 21456 31204
rect 21008 31164 21456 31192
rect 21450 31152 21456 31164
rect 21508 31152 21514 31204
rect 21910 31152 21916 31204
rect 21968 31192 21974 31204
rect 22204 31192 22232 31223
rect 21968 31164 22232 31192
rect 22296 31192 22324 31223
rect 22738 31220 22744 31272
rect 22796 31260 22802 31272
rect 22925 31263 22983 31269
rect 22925 31260 22937 31263
rect 22796 31232 22937 31260
rect 22796 31220 22802 31232
rect 22925 31229 22937 31232
rect 22971 31260 22983 31263
rect 24504 31260 24532 31291
rect 24946 31288 24952 31340
rect 25004 31328 25010 31340
rect 25593 31331 25651 31337
rect 25593 31328 25605 31331
rect 25004 31300 25605 31328
rect 25004 31288 25010 31300
rect 25593 31297 25605 31300
rect 25639 31297 25651 31331
rect 25593 31291 25651 31297
rect 25774 31288 25780 31340
rect 25832 31328 25838 31340
rect 25869 31331 25927 31337
rect 25869 31328 25881 31331
rect 25832 31300 25881 31328
rect 25832 31288 25838 31300
rect 25869 31297 25881 31300
rect 25915 31297 25927 31331
rect 25869 31291 25927 31297
rect 26145 31331 26203 31337
rect 26145 31297 26157 31331
rect 26191 31297 26203 31331
rect 26145 31291 26203 31297
rect 26329 31331 26387 31337
rect 26329 31297 26341 31331
rect 26375 31328 26387 31331
rect 26418 31328 26424 31340
rect 26375 31300 26424 31328
rect 26375 31297 26387 31300
rect 26329 31291 26387 31297
rect 22971 31232 24532 31260
rect 25961 31263 26019 31269
rect 22971 31229 22983 31232
rect 22925 31223 22983 31229
rect 25961 31229 25973 31263
rect 26007 31229 26019 31263
rect 26160 31260 26188 31291
rect 26418 31288 26424 31300
rect 26476 31328 26482 31340
rect 26786 31328 26792 31340
rect 26476 31300 26792 31328
rect 26476 31288 26482 31300
rect 26786 31288 26792 31300
rect 26844 31288 26850 31340
rect 26988 31337 27016 31368
rect 27080 31337 27108 31436
rect 27522 31424 27528 31476
rect 27580 31464 27586 31476
rect 29181 31467 29239 31473
rect 29181 31464 29193 31467
rect 27580 31436 29193 31464
rect 27580 31424 27586 31436
rect 29181 31433 29193 31436
rect 29227 31433 29239 31467
rect 29181 31427 29239 31433
rect 30558 31424 30564 31476
rect 30616 31464 30622 31476
rect 33134 31464 33140 31476
rect 30616 31436 31156 31464
rect 33095 31436 33140 31464
rect 30616 31424 30622 31436
rect 27246 31396 27252 31408
rect 27207 31368 27252 31396
rect 27246 31356 27252 31368
rect 27304 31356 27310 31408
rect 30466 31396 30472 31408
rect 28276 31368 30472 31396
rect 26973 31331 27031 31337
rect 26973 31297 26985 31331
rect 27019 31297 27031 31331
rect 26973 31291 27031 31297
rect 27066 31331 27124 31337
rect 27066 31297 27078 31331
rect 27112 31297 27124 31331
rect 27066 31291 27124 31297
rect 27264 31260 27292 31356
rect 28276 31337 28304 31368
rect 30466 31356 30472 31368
rect 30524 31356 30530 31408
rect 30668 31368 31064 31396
rect 27341 31331 27399 31337
rect 27341 31297 27353 31331
rect 27387 31297 27399 31331
rect 27341 31291 27399 31297
rect 27479 31331 27537 31337
rect 27479 31297 27491 31331
rect 27525 31328 27537 31331
rect 28261 31331 28319 31337
rect 27525 31300 28120 31328
rect 27525 31297 27537 31300
rect 27479 31291 27537 31297
rect 26160 31232 27292 31260
rect 25961 31223 26019 31229
rect 25976 31192 26004 31223
rect 26326 31192 26332 31204
rect 22296 31164 23980 31192
rect 25976 31164 26332 31192
rect 21968 31152 21974 31164
rect 23952 31136 23980 31164
rect 26326 31152 26332 31164
rect 26384 31152 26390 31204
rect 26602 31152 26608 31204
rect 26660 31192 26666 31204
rect 27356 31192 27384 31291
rect 28092 31260 28120 31300
rect 28261 31297 28273 31331
rect 28307 31297 28319 31331
rect 28261 31291 28319 31297
rect 28353 31331 28411 31337
rect 28353 31297 28365 31331
rect 28399 31328 28411 31331
rect 28534 31328 28540 31340
rect 28399 31300 28540 31328
rect 28399 31297 28411 31300
rect 28353 31291 28411 31297
rect 28534 31288 28540 31300
rect 28592 31288 28598 31340
rect 28629 31331 28687 31337
rect 28629 31297 28641 31331
rect 28675 31297 28687 31331
rect 29086 31328 29092 31340
rect 29047 31300 29092 31328
rect 28629 31291 28687 31297
rect 28092 31232 28304 31260
rect 28276 31204 28304 31232
rect 26660 31164 28212 31192
rect 26660 31152 26666 31164
rect 15286 31084 15292 31136
rect 15344 31124 15350 31136
rect 16942 31124 16948 31136
rect 15344 31096 16948 31124
rect 15344 31084 15350 31096
rect 16942 31084 16948 31096
rect 17000 31084 17006 31136
rect 18138 31124 18144 31136
rect 18099 31096 18144 31124
rect 18138 31084 18144 31096
rect 18196 31084 18202 31136
rect 19978 31084 19984 31136
rect 20036 31124 20042 31136
rect 20073 31127 20131 31133
rect 20073 31124 20085 31127
rect 20036 31096 20085 31124
rect 20036 31084 20042 31096
rect 20073 31093 20085 31096
rect 20119 31093 20131 31127
rect 20073 31087 20131 31093
rect 23198 31084 23204 31136
rect 23256 31124 23262 31136
rect 23293 31127 23351 31133
rect 23293 31124 23305 31127
rect 23256 31096 23305 31124
rect 23256 31084 23262 31096
rect 23293 31093 23305 31096
rect 23339 31093 23351 31127
rect 23934 31124 23940 31136
rect 23895 31096 23940 31124
rect 23293 31087 23351 31093
rect 23934 31084 23940 31096
rect 23992 31084 23998 31136
rect 27246 31084 27252 31136
rect 27304 31124 27310 31136
rect 27617 31127 27675 31133
rect 27617 31124 27629 31127
rect 27304 31096 27629 31124
rect 27304 31084 27310 31096
rect 27617 31093 27629 31096
rect 27663 31093 27675 31127
rect 28074 31124 28080 31136
rect 28035 31096 28080 31124
rect 27617 31087 27675 31093
rect 28074 31084 28080 31096
rect 28132 31084 28138 31136
rect 28184 31124 28212 31164
rect 28258 31152 28264 31204
rect 28316 31192 28322 31204
rect 28537 31195 28595 31201
rect 28537 31192 28549 31195
rect 28316 31164 28549 31192
rect 28316 31152 28322 31164
rect 28537 31161 28549 31164
rect 28583 31161 28595 31195
rect 28537 31155 28595 31161
rect 28644 31124 28672 31291
rect 29086 31288 29092 31300
rect 29144 31288 29150 31340
rect 29822 31288 29828 31340
rect 29880 31328 29886 31340
rect 29917 31331 29975 31337
rect 29917 31328 29929 31331
rect 29880 31300 29929 31328
rect 29880 31288 29886 31300
rect 29917 31297 29929 31300
rect 29963 31297 29975 31331
rect 29917 31291 29975 31297
rect 30561 31331 30619 31337
rect 30561 31297 30573 31331
rect 30607 31328 30619 31331
rect 30668 31328 30696 31368
rect 30607 31300 30696 31328
rect 30745 31331 30803 31337
rect 30607 31297 30619 31300
rect 30561 31291 30619 31297
rect 30745 31297 30757 31331
rect 30791 31297 30803 31331
rect 30926 31328 30932 31340
rect 30887 31300 30932 31328
rect 30745 31291 30803 31297
rect 29546 31220 29552 31272
rect 29604 31260 29610 31272
rect 29733 31263 29791 31269
rect 29733 31260 29745 31263
rect 29604 31232 29745 31260
rect 29604 31220 29610 31232
rect 29733 31229 29745 31232
rect 29779 31260 29791 31263
rect 30466 31260 30472 31272
rect 29779 31232 30472 31260
rect 29779 31229 29791 31232
rect 29733 31223 29791 31229
rect 30466 31220 30472 31232
rect 30524 31220 30530 31272
rect 29822 31152 29828 31204
rect 29880 31192 29886 31204
rect 30760 31192 30788 31291
rect 30926 31288 30932 31300
rect 30984 31288 30990 31340
rect 30837 31263 30895 31269
rect 30837 31229 30849 31263
rect 30883 31229 30895 31263
rect 31036 31260 31064 31368
rect 31128 31337 31156 31436
rect 33134 31424 33140 31436
rect 33192 31424 33198 31476
rect 31294 31356 31300 31408
rect 31352 31396 31358 31408
rect 31352 31368 33640 31396
rect 31352 31356 31358 31368
rect 31113 31331 31171 31337
rect 31113 31297 31125 31331
rect 31159 31297 31171 31331
rect 31113 31291 31171 31297
rect 31846 31288 31852 31340
rect 31904 31328 31910 31340
rect 32122 31328 32128 31340
rect 31904 31300 32128 31328
rect 31904 31288 31910 31300
rect 32122 31288 32128 31300
rect 32180 31288 32186 31340
rect 33612 31337 33640 31368
rect 32769 31331 32827 31337
rect 32769 31297 32781 31331
rect 32815 31297 32827 31331
rect 32769 31291 32827 31297
rect 33597 31331 33655 31337
rect 33597 31297 33609 31331
rect 33643 31297 33655 31331
rect 33597 31291 33655 31297
rect 33781 31331 33839 31337
rect 33781 31297 33793 31331
rect 33827 31297 33839 31331
rect 34514 31328 34520 31340
rect 34475 31300 34520 31328
rect 33781 31291 33839 31297
rect 32030 31260 32036 31272
rect 31036 31232 32036 31260
rect 30837 31223 30895 31229
rect 29880 31164 30788 31192
rect 29880 31152 29886 31164
rect 30098 31124 30104 31136
rect 28184 31096 28672 31124
rect 30059 31096 30104 31124
rect 30098 31084 30104 31096
rect 30156 31084 30162 31136
rect 30466 31084 30472 31136
rect 30524 31124 30530 31136
rect 30852 31124 30880 31223
rect 32030 31220 32036 31232
rect 32088 31220 32094 31272
rect 32582 31220 32588 31272
rect 32640 31260 32646 31272
rect 32677 31263 32735 31269
rect 32677 31260 32689 31263
rect 32640 31232 32689 31260
rect 32640 31220 32646 31232
rect 32677 31229 32689 31232
rect 32723 31229 32735 31263
rect 32784 31260 32812 31291
rect 32858 31260 32864 31272
rect 32784 31232 32864 31260
rect 32677 31223 32735 31229
rect 32858 31220 32864 31232
rect 32916 31260 32922 31272
rect 33796 31260 33824 31291
rect 34514 31288 34520 31300
rect 34572 31288 34578 31340
rect 35526 31328 35532 31340
rect 35487 31300 35532 31328
rect 35526 31288 35532 31300
rect 35584 31288 35590 31340
rect 34606 31260 34612 31272
rect 32916 31232 33824 31260
rect 34567 31232 34612 31260
rect 32916 31220 32922 31232
rect 34606 31220 34612 31232
rect 34664 31220 34670 31272
rect 34885 31263 34943 31269
rect 34885 31229 34897 31263
rect 34931 31260 34943 31263
rect 35437 31263 35495 31269
rect 35437 31260 35449 31263
rect 34931 31232 35449 31260
rect 34931 31229 34943 31232
rect 34885 31223 34943 31229
rect 35437 31229 35449 31232
rect 35483 31229 35495 31263
rect 35437 31223 35495 31229
rect 31202 31152 31208 31204
rect 31260 31192 31266 31204
rect 33597 31195 33655 31201
rect 33597 31192 33609 31195
rect 31260 31164 33609 31192
rect 31260 31152 31266 31164
rect 33597 31161 33609 31164
rect 33643 31161 33655 31195
rect 33597 31155 33655 31161
rect 35897 31195 35955 31201
rect 35897 31161 35909 31195
rect 35943 31192 35955 31195
rect 35986 31192 35992 31204
rect 35943 31164 35992 31192
rect 35943 31161 35955 31164
rect 35897 31155 35955 31161
rect 35986 31152 35992 31164
rect 36044 31152 36050 31204
rect 30524 31096 30880 31124
rect 31297 31127 31355 31133
rect 30524 31084 30530 31096
rect 31297 31093 31309 31127
rect 31343 31124 31355 31127
rect 31478 31124 31484 31136
rect 31343 31096 31484 31124
rect 31343 31093 31355 31096
rect 31297 31087 31355 31093
rect 31478 31084 31484 31096
rect 31536 31084 31542 31136
rect 31662 31084 31668 31136
rect 31720 31124 31726 31136
rect 32674 31124 32680 31136
rect 31720 31096 32680 31124
rect 31720 31084 31726 31096
rect 32674 31084 32680 31096
rect 32732 31084 32738 31136
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 15194 30920 15200 30932
rect 15155 30892 15200 30920
rect 15194 30880 15200 30892
rect 15252 30880 15258 30932
rect 16393 30923 16451 30929
rect 16393 30889 16405 30923
rect 16439 30920 16451 30923
rect 16758 30920 16764 30932
rect 16439 30892 16764 30920
rect 16439 30889 16451 30892
rect 16393 30883 16451 30889
rect 16758 30880 16764 30892
rect 16816 30880 16822 30932
rect 18230 30920 18236 30932
rect 17788 30892 18236 30920
rect 16022 30784 16028 30796
rect 15580 30756 16028 30784
rect 15580 30725 15608 30756
rect 16022 30744 16028 30756
rect 16080 30744 16086 30796
rect 15473 30719 15531 30725
rect 15473 30685 15485 30719
rect 15519 30685 15531 30719
rect 15473 30679 15531 30685
rect 15565 30719 15623 30725
rect 15565 30685 15577 30719
rect 15611 30685 15623 30719
rect 15565 30679 15623 30685
rect 15488 30648 15516 30679
rect 15654 30676 15660 30728
rect 15712 30716 15718 30728
rect 15841 30719 15899 30725
rect 15712 30688 15757 30716
rect 15712 30676 15718 30688
rect 15841 30685 15853 30719
rect 15887 30716 15899 30719
rect 15930 30716 15936 30728
rect 15887 30688 15936 30716
rect 15887 30685 15899 30688
rect 15841 30679 15899 30685
rect 15930 30676 15936 30688
rect 15988 30676 15994 30728
rect 16574 30716 16580 30728
rect 16535 30688 16580 30716
rect 16574 30676 16580 30688
rect 16632 30676 16638 30728
rect 16853 30719 16911 30725
rect 16853 30685 16865 30719
rect 16899 30716 16911 30719
rect 17037 30719 17095 30725
rect 16899 30688 16988 30716
rect 16899 30685 16911 30688
rect 16853 30679 16911 30685
rect 16669 30651 16727 30657
rect 15488 30620 15884 30648
rect 15856 30592 15884 30620
rect 16669 30617 16681 30651
rect 16715 30617 16727 30651
rect 16669 30611 16727 30617
rect 15838 30540 15844 30592
rect 15896 30540 15902 30592
rect 16684 30580 16712 30611
rect 16758 30608 16764 30660
rect 16816 30648 16822 30660
rect 16960 30648 16988 30688
rect 17037 30685 17049 30719
rect 17083 30716 17095 30719
rect 17586 30716 17592 30728
rect 17083 30688 17592 30716
rect 17083 30685 17095 30688
rect 17037 30679 17095 30685
rect 17586 30676 17592 30688
rect 17644 30676 17650 30728
rect 17788 30725 17816 30892
rect 18230 30880 18236 30892
rect 18288 30880 18294 30932
rect 20070 30880 20076 30932
rect 20128 30920 20134 30932
rect 20717 30923 20775 30929
rect 20717 30920 20729 30923
rect 20128 30892 20729 30920
rect 20128 30880 20134 30892
rect 20717 30889 20729 30892
rect 20763 30889 20775 30923
rect 20717 30883 20775 30889
rect 21082 30880 21088 30932
rect 21140 30920 21146 30932
rect 21269 30923 21327 30929
rect 21269 30920 21281 30923
rect 21140 30892 21281 30920
rect 21140 30880 21146 30892
rect 21269 30889 21281 30892
rect 21315 30889 21327 30923
rect 21269 30883 21327 30889
rect 23106 30880 23112 30932
rect 23164 30920 23170 30932
rect 29730 30920 29736 30932
rect 23164 30892 29040 30920
rect 29691 30892 29736 30920
rect 23164 30880 23170 30892
rect 17954 30812 17960 30864
rect 18012 30812 18018 30864
rect 18138 30852 18144 30864
rect 18099 30824 18144 30852
rect 18138 30812 18144 30824
rect 18196 30812 18202 30864
rect 19245 30855 19303 30861
rect 19245 30821 19257 30855
rect 19291 30852 19303 30855
rect 23014 30852 23020 30864
rect 19291 30824 23020 30852
rect 19291 30821 19303 30824
rect 19245 30815 19303 30821
rect 23014 30812 23020 30824
rect 23072 30812 23078 30864
rect 23474 30852 23480 30864
rect 23435 30824 23480 30852
rect 23474 30812 23480 30824
rect 23532 30812 23538 30864
rect 24946 30812 24952 30864
rect 25004 30852 25010 30864
rect 25225 30855 25283 30861
rect 25225 30852 25237 30855
rect 25004 30824 25237 30852
rect 25004 30812 25010 30824
rect 25225 30821 25237 30824
rect 25271 30821 25283 30855
rect 28902 30852 28908 30864
rect 25225 30815 25283 30821
rect 26896 30824 28908 30852
rect 17972 30725 18000 30812
rect 18156 30784 18184 30812
rect 23198 30784 23204 30796
rect 18156 30756 21772 30784
rect 23159 30756 23204 30784
rect 17773 30719 17831 30725
rect 17773 30685 17785 30719
rect 17819 30685 17831 30719
rect 17957 30719 18015 30725
rect 17957 30716 17969 30719
rect 17773 30679 17831 30685
rect 17880 30688 17969 30716
rect 16816 30620 16861 30648
rect 16960 30620 17816 30648
rect 16816 30608 16822 30620
rect 17788 30592 17816 30620
rect 17034 30580 17040 30592
rect 16684 30552 17040 30580
rect 17034 30540 17040 30552
rect 17092 30540 17098 30592
rect 17770 30540 17776 30592
rect 17828 30540 17834 30592
rect 17880 30580 17908 30688
rect 17957 30685 17969 30688
rect 18003 30685 18015 30719
rect 17957 30679 18015 30685
rect 18046 30676 18052 30728
rect 18104 30716 18110 30728
rect 18141 30719 18199 30725
rect 18141 30716 18153 30719
rect 18104 30688 18153 30716
rect 18104 30676 18110 30688
rect 18141 30685 18153 30688
rect 18187 30685 18199 30719
rect 18141 30679 18199 30685
rect 18322 30676 18328 30728
rect 18380 30716 18386 30728
rect 18509 30719 18567 30725
rect 18509 30716 18521 30719
rect 18380 30688 18521 30716
rect 18380 30676 18386 30688
rect 18509 30685 18521 30688
rect 18555 30716 18567 30719
rect 19429 30719 19487 30725
rect 19429 30716 19441 30719
rect 18555 30688 19441 30716
rect 18555 30685 18567 30688
rect 18509 30679 18567 30685
rect 19429 30685 19441 30688
rect 19475 30716 19487 30719
rect 19518 30716 19524 30728
rect 19475 30688 19524 30716
rect 19475 30685 19487 30688
rect 19429 30679 19487 30685
rect 19518 30676 19524 30688
rect 19576 30676 19582 30728
rect 19705 30719 19763 30725
rect 19705 30716 19717 30719
rect 19628 30688 19717 30716
rect 19334 30608 19340 30660
rect 19392 30648 19398 30660
rect 19628 30648 19656 30688
rect 19705 30685 19717 30688
rect 19751 30685 19763 30719
rect 19705 30679 19763 30685
rect 20441 30719 20499 30725
rect 20441 30685 20453 30719
rect 20487 30685 20499 30719
rect 20441 30679 20499 30685
rect 20533 30719 20591 30725
rect 20533 30685 20545 30719
rect 20579 30716 20591 30719
rect 21450 30716 21456 30728
rect 20579 30688 21456 30716
rect 20579 30685 20591 30688
rect 20533 30679 20591 30685
rect 19392 30620 19656 30648
rect 20456 30648 20484 30679
rect 21450 30676 21456 30688
rect 21508 30676 21514 30728
rect 21744 30725 21772 30756
rect 23198 30744 23204 30756
rect 23256 30744 23262 30796
rect 26694 30784 26700 30796
rect 26068 30756 26700 30784
rect 21729 30719 21787 30725
rect 21729 30685 21741 30719
rect 21775 30716 21787 30719
rect 22186 30716 22192 30728
rect 21775 30688 22094 30716
rect 22147 30688 22192 30716
rect 21775 30685 21787 30688
rect 21729 30679 21787 30685
rect 21266 30648 21272 30660
rect 20456 30620 21272 30648
rect 19392 30608 19398 30620
rect 21266 30608 21272 30620
rect 21324 30608 21330 30660
rect 22066 30648 22094 30688
rect 22186 30676 22192 30688
rect 22244 30676 22250 30728
rect 22370 30716 22376 30728
rect 22331 30688 22376 30716
rect 22370 30676 22376 30688
rect 22428 30676 22434 30728
rect 23109 30719 23167 30725
rect 23109 30685 23121 30719
rect 23155 30716 23167 30719
rect 23934 30716 23940 30728
rect 23155 30688 23940 30716
rect 23155 30685 23167 30688
rect 23109 30679 23167 30685
rect 23934 30676 23940 30688
rect 23992 30676 23998 30728
rect 26068 30725 26096 30756
rect 26694 30744 26700 30756
rect 26752 30744 26758 30796
rect 26053 30719 26111 30725
rect 26053 30685 26065 30719
rect 26099 30685 26111 30719
rect 26234 30716 26240 30728
rect 26195 30688 26240 30716
rect 26053 30679 26111 30685
rect 26234 30676 26240 30688
rect 26292 30676 26298 30728
rect 26896 30725 26924 30824
rect 28902 30812 28908 30824
rect 28960 30812 28966 30864
rect 28074 30784 28080 30796
rect 26988 30756 28080 30784
rect 26988 30725 27016 30756
rect 28074 30744 28080 30756
rect 28132 30744 28138 30796
rect 28261 30787 28319 30793
rect 28261 30753 28273 30787
rect 28307 30784 28319 30787
rect 28350 30784 28356 30796
rect 28307 30756 28356 30784
rect 28307 30753 28319 30756
rect 28261 30747 28319 30753
rect 28350 30744 28356 30756
rect 28408 30744 28414 30796
rect 29012 30784 29040 30892
rect 29730 30880 29736 30892
rect 29788 30880 29794 30932
rect 30374 30880 30380 30932
rect 30432 30920 30438 30932
rect 30653 30923 30711 30929
rect 30653 30920 30665 30923
rect 30432 30892 30665 30920
rect 30432 30880 30438 30892
rect 30653 30889 30665 30892
rect 30699 30889 30711 30923
rect 30653 30883 30711 30889
rect 31018 30880 31024 30932
rect 31076 30920 31082 30932
rect 31113 30923 31171 30929
rect 31113 30920 31125 30923
rect 31076 30892 31125 30920
rect 31076 30880 31082 30892
rect 31113 30889 31125 30892
rect 31159 30889 31171 30923
rect 31478 30920 31484 30932
rect 31439 30892 31484 30920
rect 31113 30883 31171 30889
rect 31478 30880 31484 30892
rect 31536 30880 31542 30932
rect 31570 30880 31576 30932
rect 31628 30920 31634 30932
rect 32493 30923 32551 30929
rect 31628 30892 31673 30920
rect 31628 30880 31634 30892
rect 32493 30889 32505 30923
rect 32539 30889 32551 30923
rect 32674 30920 32680 30932
rect 32635 30892 32680 30920
rect 32493 30883 32551 30889
rect 30098 30812 30104 30864
rect 30156 30852 30162 30864
rect 31389 30855 31447 30861
rect 31389 30852 31401 30855
rect 30156 30824 31401 30852
rect 30156 30812 30162 30824
rect 31389 30821 31401 30824
rect 31435 30821 31447 30855
rect 31846 30852 31852 30864
rect 31389 30815 31447 30821
rect 31496 30824 31852 30852
rect 31496 30784 31524 30824
rect 31846 30812 31852 30824
rect 31904 30812 31910 30864
rect 32508 30852 32536 30883
rect 32674 30880 32680 30892
rect 32732 30880 32738 30932
rect 33413 30923 33471 30929
rect 33413 30889 33425 30923
rect 33459 30920 33471 30923
rect 33962 30920 33968 30932
rect 33459 30892 33968 30920
rect 33459 30889 33471 30892
rect 33413 30883 33471 30889
rect 33962 30880 33968 30892
rect 34020 30880 34026 30932
rect 33318 30852 33324 30864
rect 32508 30824 33324 30852
rect 29012 30756 31524 30784
rect 31570 30744 31576 30796
rect 31628 30784 31634 30796
rect 32508 30784 32536 30824
rect 33318 30812 33324 30824
rect 33376 30812 33382 30864
rect 35986 30784 35992 30796
rect 31628 30756 31800 30784
rect 31628 30744 31634 30756
rect 26881 30719 26939 30725
rect 26881 30685 26893 30719
rect 26927 30685 26939 30719
rect 26881 30679 26939 30685
rect 26973 30719 27031 30725
rect 26973 30685 26985 30719
rect 27019 30685 27031 30719
rect 26973 30679 27031 30685
rect 27157 30719 27215 30725
rect 27157 30685 27169 30719
rect 27203 30685 27215 30719
rect 27157 30679 27215 30685
rect 22830 30648 22836 30660
rect 22066 30620 22836 30648
rect 22830 30608 22836 30620
rect 22888 30608 22894 30660
rect 24949 30651 25007 30657
rect 24949 30617 24961 30651
rect 24995 30648 25007 30651
rect 25222 30648 25228 30660
rect 24995 30620 25228 30648
rect 24995 30617 25007 30620
rect 24949 30611 25007 30617
rect 25222 30608 25228 30620
rect 25280 30608 25286 30660
rect 26326 30608 26332 30660
rect 26384 30648 26390 30660
rect 27172 30648 27200 30679
rect 27246 30676 27252 30728
rect 27304 30716 27310 30728
rect 28169 30719 28227 30725
rect 27304 30688 27349 30716
rect 27304 30676 27310 30688
rect 28169 30685 28181 30719
rect 28215 30716 28227 30719
rect 28534 30716 28540 30728
rect 28215 30688 28540 30716
rect 28215 30685 28227 30688
rect 28169 30679 28227 30685
rect 28534 30676 28540 30688
rect 28592 30676 28598 30728
rect 28721 30719 28779 30725
rect 28721 30685 28733 30719
rect 28767 30716 28779 30719
rect 28994 30716 29000 30728
rect 28767 30688 29000 30716
rect 28767 30685 28779 30688
rect 28721 30679 28779 30685
rect 28994 30676 29000 30688
rect 29052 30676 29058 30728
rect 30285 30719 30343 30725
rect 30285 30685 30297 30719
rect 30331 30716 30343 30719
rect 31110 30716 31116 30728
rect 30331 30688 31116 30716
rect 30331 30685 30343 30688
rect 30285 30679 30343 30685
rect 31110 30676 31116 30688
rect 31168 30676 31174 30728
rect 31665 30719 31723 30725
rect 31665 30685 31677 30719
rect 31711 30685 31723 30719
rect 31665 30679 31723 30685
rect 26384 30620 27200 30648
rect 29641 30651 29699 30657
rect 26384 30608 26390 30620
rect 29641 30617 29653 30651
rect 29687 30648 29699 30651
rect 30469 30651 30527 30657
rect 29687 30620 30328 30648
rect 29687 30617 29699 30620
rect 29641 30611 29699 30617
rect 30300 30592 30328 30620
rect 30469 30617 30481 30651
rect 30515 30648 30527 30651
rect 30926 30648 30932 30660
rect 30515 30620 30932 30648
rect 30515 30617 30527 30620
rect 30469 30611 30527 30617
rect 30926 30608 30932 30620
rect 30984 30648 30990 30660
rect 31386 30648 31392 30660
rect 30984 30620 31392 30648
rect 30984 30608 30990 30620
rect 31386 30608 31392 30620
rect 31444 30608 31450 30660
rect 18046 30580 18052 30592
rect 17880 30552 18052 30580
rect 18046 30540 18052 30552
rect 18104 30540 18110 30592
rect 18598 30540 18604 30592
rect 18656 30580 18662 30592
rect 19613 30583 19671 30589
rect 19613 30580 19625 30583
rect 18656 30552 19625 30580
rect 18656 30540 18662 30552
rect 19613 30549 19625 30552
rect 19659 30580 19671 30583
rect 21634 30580 21640 30592
rect 19659 30552 21640 30580
rect 19659 30549 19671 30552
rect 19613 30543 19671 30549
rect 21634 30540 21640 30552
rect 21692 30540 21698 30592
rect 21726 30540 21732 30592
rect 21784 30580 21790 30592
rect 22281 30583 22339 30589
rect 22281 30580 22293 30583
rect 21784 30552 22293 30580
rect 21784 30540 21790 30552
rect 22281 30549 22293 30552
rect 22327 30549 22339 30583
rect 25406 30580 25412 30592
rect 25367 30552 25412 30580
rect 22281 30543 22339 30549
rect 25406 30540 25412 30552
rect 25464 30540 25470 30592
rect 26142 30580 26148 30592
rect 26103 30552 26148 30580
rect 26142 30540 26148 30552
rect 26200 30540 26206 30592
rect 26697 30583 26755 30589
rect 26697 30549 26709 30583
rect 26743 30580 26755 30583
rect 27338 30580 27344 30592
rect 26743 30552 27344 30580
rect 26743 30549 26755 30552
rect 26697 30543 26755 30549
rect 27338 30540 27344 30552
rect 27396 30540 27402 30592
rect 28810 30540 28816 30592
rect 28868 30580 28874 30592
rect 28905 30583 28963 30589
rect 28905 30580 28917 30583
rect 28868 30552 28917 30580
rect 28868 30540 28874 30552
rect 28905 30549 28917 30552
rect 28951 30580 28963 30583
rect 29454 30580 29460 30592
rect 28951 30552 29460 30580
rect 28951 30549 28963 30552
rect 28905 30543 28963 30549
rect 29454 30540 29460 30552
rect 29512 30540 29518 30592
rect 30282 30540 30288 30592
rect 30340 30540 30346 30592
rect 31680 30580 31708 30679
rect 31772 30648 31800 30756
rect 31864 30756 32536 30784
rect 35947 30756 35992 30784
rect 31864 30725 31892 30756
rect 35986 30744 35992 30756
rect 36044 30744 36050 30796
rect 31849 30719 31907 30725
rect 31849 30685 31861 30719
rect 31895 30685 31907 30719
rect 31849 30679 31907 30685
rect 32309 30719 32367 30725
rect 32309 30685 32321 30719
rect 32355 30685 32367 30719
rect 32309 30679 32367 30685
rect 32493 30719 32551 30725
rect 32493 30685 32505 30719
rect 32539 30685 32551 30719
rect 32493 30679 32551 30685
rect 32324 30648 32352 30679
rect 31772 30620 32352 30648
rect 32508 30648 32536 30679
rect 32582 30676 32588 30728
rect 32640 30716 32646 30728
rect 33413 30719 33471 30725
rect 33413 30716 33425 30719
rect 32640 30688 33425 30716
rect 32640 30676 32646 30688
rect 33413 30685 33425 30688
rect 33459 30685 33471 30719
rect 33594 30716 33600 30728
rect 33555 30688 33600 30716
rect 33413 30679 33471 30685
rect 32766 30648 32772 30660
rect 32508 30620 32772 30648
rect 32122 30580 32128 30592
rect 31680 30552 32128 30580
rect 32122 30540 32128 30552
rect 32180 30580 32186 30592
rect 32508 30580 32536 30620
rect 32766 30608 32772 30620
rect 32824 30608 32830 30660
rect 33428 30648 33456 30679
rect 33594 30676 33600 30688
rect 33652 30676 33658 30728
rect 35066 30716 35072 30728
rect 35027 30688 35072 30716
rect 35066 30676 35072 30688
rect 35124 30676 35130 30728
rect 35253 30719 35311 30725
rect 35253 30685 35265 30719
rect 35299 30716 35311 30719
rect 35618 30716 35624 30728
rect 35299 30688 35624 30716
rect 35299 30685 35311 30688
rect 35253 30679 35311 30685
rect 35618 30676 35624 30688
rect 35676 30676 35682 30728
rect 35894 30716 35900 30728
rect 35855 30688 35900 30716
rect 35894 30676 35900 30688
rect 35952 30676 35958 30728
rect 34054 30648 34060 30660
rect 33428 30620 34060 30648
rect 34054 30608 34060 30620
rect 34112 30608 34118 30660
rect 32180 30552 32536 30580
rect 35161 30583 35219 30589
rect 32180 30540 32186 30552
rect 35161 30549 35173 30583
rect 35207 30580 35219 30583
rect 36170 30580 36176 30592
rect 35207 30552 36176 30580
rect 35207 30549 35219 30552
rect 35161 30543 35219 30549
rect 36170 30540 36176 30552
rect 36228 30540 36234 30592
rect 36265 30583 36323 30589
rect 36265 30549 36277 30583
rect 36311 30580 36323 30583
rect 37182 30580 37188 30592
rect 36311 30552 37188 30580
rect 36311 30549 36323 30552
rect 36265 30543 36323 30549
rect 37182 30540 37188 30552
rect 37240 30540 37246 30592
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 15930 30376 15936 30388
rect 15580 30348 15936 30376
rect 15580 30249 15608 30348
rect 15654 30268 15660 30320
rect 15712 30308 15718 30320
rect 15749 30311 15807 30317
rect 15749 30308 15761 30311
rect 15712 30280 15761 30308
rect 15712 30268 15718 30280
rect 15749 30277 15761 30280
rect 15795 30277 15807 30311
rect 15856 30308 15884 30348
rect 15930 30336 15936 30348
rect 15988 30336 15994 30388
rect 17862 30336 17868 30388
rect 17920 30376 17926 30388
rect 18322 30376 18328 30388
rect 17920 30348 18328 30376
rect 17920 30336 17926 30348
rect 18322 30336 18328 30348
rect 18380 30336 18386 30388
rect 18506 30376 18512 30388
rect 18467 30348 18512 30376
rect 18506 30336 18512 30348
rect 18564 30336 18570 30388
rect 18969 30379 19027 30385
rect 18969 30345 18981 30379
rect 19015 30345 19027 30379
rect 18969 30339 19027 30345
rect 18984 30308 19012 30339
rect 21450 30336 21456 30388
rect 21508 30376 21514 30388
rect 22094 30376 22100 30388
rect 21508 30348 22100 30376
rect 21508 30336 21514 30348
rect 22094 30336 22100 30348
rect 22152 30336 22158 30388
rect 22189 30379 22247 30385
rect 22189 30345 22201 30379
rect 22235 30376 22247 30379
rect 22738 30376 22744 30388
rect 22235 30348 22744 30376
rect 22235 30345 22247 30348
rect 22189 30339 22247 30345
rect 22738 30336 22744 30348
rect 22796 30336 22802 30388
rect 22859 30379 22917 30385
rect 22859 30345 22871 30379
rect 22905 30376 22917 30379
rect 23198 30376 23204 30388
rect 22905 30348 23204 30376
rect 22905 30345 22917 30348
rect 22859 30339 22917 30345
rect 23198 30336 23204 30348
rect 23256 30376 23262 30388
rect 23842 30376 23848 30388
rect 23256 30348 23848 30376
rect 23256 30336 23262 30348
rect 23842 30336 23848 30348
rect 23900 30336 23906 30388
rect 26234 30336 26240 30388
rect 26292 30376 26298 30388
rect 28534 30376 28540 30388
rect 26292 30348 28540 30376
rect 26292 30336 26298 30348
rect 28534 30336 28540 30348
rect 28592 30336 28598 30388
rect 30374 30336 30380 30388
rect 30432 30376 30438 30388
rect 31294 30376 31300 30388
rect 30432 30348 31300 30376
rect 30432 30336 30438 30348
rect 31294 30336 31300 30348
rect 31352 30336 31358 30388
rect 34885 30379 34943 30385
rect 34885 30345 34897 30379
rect 34931 30376 34943 30379
rect 35066 30376 35072 30388
rect 34931 30348 35072 30376
rect 34931 30345 34943 30348
rect 34885 30339 34943 30345
rect 35066 30336 35072 30348
rect 35124 30336 35130 30388
rect 20806 30308 20812 30320
rect 15856 30280 19012 30308
rect 20767 30280 20812 30308
rect 15749 30271 15807 30277
rect 20806 30268 20812 30280
rect 20864 30268 20870 30320
rect 21634 30268 21640 30320
rect 21692 30308 21698 30320
rect 22649 30311 22707 30317
rect 22649 30308 22661 30311
rect 21692 30280 22661 30308
rect 21692 30268 21698 30280
rect 22649 30277 22661 30280
rect 22695 30277 22707 30311
rect 22649 30271 22707 30277
rect 23753 30311 23811 30317
rect 23753 30277 23765 30311
rect 23799 30308 23811 30311
rect 24118 30308 24124 30320
rect 23799 30280 24124 30308
rect 23799 30277 23811 30280
rect 23753 30271 23811 30277
rect 24118 30268 24124 30280
rect 24176 30268 24182 30320
rect 27709 30311 27767 30317
rect 27709 30308 27721 30311
rect 27540 30280 27721 30308
rect 15565 30243 15623 30249
rect 15565 30209 15577 30243
rect 15611 30209 15623 30243
rect 15838 30240 15844 30252
rect 15799 30212 15844 30240
rect 15565 30203 15623 30209
rect 15838 30200 15844 30212
rect 15896 30200 15902 30252
rect 15933 30243 15991 30249
rect 15933 30209 15945 30243
rect 15979 30240 15991 30243
rect 16574 30240 16580 30252
rect 15979 30212 16068 30240
rect 15979 30209 15991 30212
rect 15933 30203 15991 30209
rect 16040 30036 16068 30212
rect 16132 30212 16580 30240
rect 16132 30113 16160 30212
rect 16574 30200 16580 30212
rect 16632 30240 16638 30252
rect 16669 30243 16727 30249
rect 16669 30240 16681 30243
rect 16632 30212 16681 30240
rect 16632 30200 16638 30212
rect 16669 30209 16681 30212
rect 16715 30209 16727 30243
rect 17034 30240 17040 30252
rect 16995 30212 17040 30240
rect 16669 30203 16727 30209
rect 17034 30200 17040 30212
rect 17092 30200 17098 30252
rect 17405 30243 17463 30249
rect 17405 30209 17417 30243
rect 17451 30209 17463 30243
rect 17405 30203 17463 30209
rect 16758 30132 16764 30184
rect 16816 30172 16822 30184
rect 17420 30172 17448 30203
rect 17586 30200 17592 30252
rect 17644 30240 17650 30252
rect 18233 30243 18291 30249
rect 18233 30240 18245 30243
rect 17644 30212 18245 30240
rect 17644 30200 17650 30212
rect 18233 30209 18245 30212
rect 18279 30209 18291 30243
rect 19242 30240 19248 30252
rect 19203 30212 19248 30240
rect 18233 30203 18291 30209
rect 19242 30200 19248 30212
rect 19300 30200 19306 30252
rect 19426 30240 19432 30252
rect 19387 30212 19432 30240
rect 19426 30200 19432 30212
rect 19484 30200 19490 30252
rect 20073 30243 20131 30249
rect 20073 30209 20085 30243
rect 20119 30240 20131 30243
rect 20346 30240 20352 30252
rect 20119 30212 20352 30240
rect 20119 30209 20131 30212
rect 20073 30203 20131 30209
rect 17770 30172 17776 30184
rect 16816 30144 17448 30172
rect 17731 30144 17776 30172
rect 16816 30132 16822 30144
rect 17770 30132 17776 30144
rect 17828 30132 17834 30184
rect 19150 30172 19156 30184
rect 19111 30144 19156 30172
rect 19150 30132 19156 30144
rect 19208 30132 19214 30184
rect 19337 30175 19395 30181
rect 19337 30141 19349 30175
rect 19383 30172 19395 30175
rect 20088 30172 20116 30203
rect 20346 30200 20352 30212
rect 20404 30200 20410 30252
rect 20717 30243 20775 30249
rect 20717 30209 20729 30243
rect 20763 30240 20775 30243
rect 21358 30240 21364 30252
rect 20763 30212 21364 30240
rect 20763 30209 20775 30212
rect 20717 30203 20775 30209
rect 21358 30200 21364 30212
rect 21416 30200 21422 30252
rect 21818 30240 21824 30252
rect 21779 30212 21824 30240
rect 21818 30200 21824 30212
rect 21876 30200 21882 30252
rect 22002 30240 22008 30252
rect 21963 30212 22008 30240
rect 22002 30200 22008 30212
rect 22060 30200 22066 30252
rect 22738 30200 22744 30252
rect 22796 30240 22802 30252
rect 23569 30243 23627 30249
rect 23569 30240 23581 30243
rect 22796 30212 23581 30240
rect 22796 30200 22802 30212
rect 23569 30209 23581 30212
rect 23615 30209 23627 30243
rect 23569 30203 23627 30209
rect 24489 30243 24547 30249
rect 24489 30209 24501 30243
rect 24535 30240 24547 30243
rect 24578 30240 24584 30252
rect 24535 30212 24584 30240
rect 24535 30209 24547 30212
rect 24489 30203 24547 30209
rect 24578 30200 24584 30212
rect 24636 30200 24642 30252
rect 25222 30240 25228 30252
rect 25183 30212 25228 30240
rect 25222 30200 25228 30212
rect 25280 30200 25286 30252
rect 25314 30200 25320 30252
rect 25372 30240 25378 30252
rect 25869 30243 25927 30249
rect 25869 30240 25881 30243
rect 25372 30212 25881 30240
rect 25372 30200 25378 30212
rect 25869 30209 25881 30212
rect 25915 30240 25927 30243
rect 26142 30240 26148 30252
rect 25915 30212 26148 30240
rect 25915 30209 25927 30212
rect 25869 30203 25927 30209
rect 26142 30200 26148 30212
rect 26200 30200 26206 30252
rect 26510 30200 26516 30252
rect 26568 30240 26574 30252
rect 27540 30240 27568 30280
rect 27709 30277 27721 30280
rect 27755 30277 27767 30311
rect 27709 30271 27767 30277
rect 28074 30268 28080 30320
rect 28132 30308 28138 30320
rect 29086 30308 29092 30320
rect 28132 30280 29092 30308
rect 28132 30268 28138 30280
rect 29086 30268 29092 30280
rect 29144 30268 29150 30320
rect 29840 30280 32168 30308
rect 26568 30212 27568 30240
rect 27617 30243 27675 30249
rect 27617 30218 27629 30243
rect 27663 30218 27675 30243
rect 26568 30200 26574 30212
rect 20254 30172 20260 30184
rect 19383 30144 20116 30172
rect 20167 30144 20260 30172
rect 19383 30141 19395 30144
rect 19337 30135 19395 30141
rect 20254 30132 20260 30144
rect 20312 30172 20318 30184
rect 23106 30172 23112 30184
rect 20312 30144 23112 30172
rect 20312 30132 20318 30144
rect 23106 30132 23112 30144
rect 23164 30132 23170 30184
rect 24305 30175 24363 30181
rect 24305 30141 24317 30175
rect 24351 30172 24363 30175
rect 25038 30172 25044 30184
rect 24351 30144 25044 30172
rect 24351 30141 24363 30144
rect 24305 30135 24363 30141
rect 25038 30132 25044 30144
rect 25096 30132 25102 30184
rect 25961 30175 26019 30181
rect 25961 30172 25973 30175
rect 25332 30144 25973 30172
rect 16117 30107 16175 30113
rect 16117 30073 16129 30107
rect 16163 30073 16175 30107
rect 16117 30067 16175 30073
rect 16942 30064 16948 30116
rect 17000 30104 17006 30116
rect 22462 30104 22468 30116
rect 17000 30076 22468 30104
rect 17000 30064 17006 30076
rect 22462 30064 22468 30076
rect 22520 30064 22526 30116
rect 23566 30104 23572 30116
rect 22664 30076 23572 30104
rect 22664 30048 22692 30076
rect 23566 30064 23572 30076
rect 23624 30064 23630 30116
rect 24118 30064 24124 30116
rect 24176 30104 24182 30116
rect 24762 30104 24768 30116
rect 24176 30076 24768 30104
rect 24176 30064 24182 30076
rect 24762 30064 24768 30076
rect 24820 30064 24826 30116
rect 24946 30064 24952 30116
rect 25004 30104 25010 30116
rect 25332 30104 25360 30144
rect 25961 30141 25973 30144
rect 26007 30141 26019 30175
rect 27522 30172 27528 30184
rect 25961 30135 26019 30141
rect 26436 30144 27528 30172
rect 25004 30076 25360 30104
rect 25409 30107 25467 30113
rect 25004 30064 25010 30076
rect 25409 30073 25421 30107
rect 25455 30104 25467 30107
rect 26436 30104 26464 30144
rect 27522 30132 27528 30144
rect 27580 30132 27586 30184
rect 27614 30166 27620 30218
rect 27672 30166 27678 30218
rect 27798 30200 27804 30252
rect 27856 30240 27862 30252
rect 27939 30243 27997 30249
rect 27856 30212 27901 30240
rect 27856 30200 27862 30212
rect 27939 30209 27951 30243
rect 27985 30240 27997 30243
rect 28442 30240 28448 30252
rect 27985 30212 28448 30240
rect 27985 30209 27997 30212
rect 27939 30203 27997 30209
rect 28442 30200 28448 30212
rect 28500 30200 28506 30252
rect 28721 30243 28779 30249
rect 28721 30209 28733 30243
rect 28767 30240 28779 30243
rect 29730 30240 29736 30252
rect 28767 30212 29736 30240
rect 28767 30209 28779 30212
rect 28721 30203 28779 30209
rect 29730 30200 29736 30212
rect 29788 30200 29794 30252
rect 28077 30175 28135 30181
rect 28077 30141 28089 30175
rect 28123 30172 28135 30175
rect 28166 30172 28172 30184
rect 28123 30144 28172 30172
rect 28123 30141 28135 30144
rect 28077 30135 28135 30141
rect 28166 30132 28172 30144
rect 28224 30132 28230 30184
rect 28258 30132 28264 30184
rect 28316 30172 28322 30184
rect 29840 30172 29868 30280
rect 31389 30243 31447 30249
rect 31389 30209 31401 30243
rect 31435 30240 31447 30243
rect 31938 30240 31944 30252
rect 31435 30212 31944 30240
rect 31435 30209 31447 30212
rect 31389 30203 31447 30209
rect 31938 30200 31944 30212
rect 31996 30200 32002 30252
rect 32140 30249 32168 30280
rect 32214 30268 32220 30320
rect 32272 30308 32278 30320
rect 32309 30311 32367 30317
rect 32309 30308 32321 30311
rect 32272 30280 32321 30308
rect 32272 30268 32278 30280
rect 32309 30277 32321 30280
rect 32355 30277 32367 30311
rect 32950 30308 32956 30320
rect 32309 30271 32367 30277
rect 32416 30280 32956 30308
rect 32416 30249 32444 30280
rect 32950 30268 32956 30280
rect 33008 30268 33014 30320
rect 33965 30311 34023 30317
rect 33965 30277 33977 30311
rect 34011 30308 34023 30311
rect 35618 30308 35624 30320
rect 34011 30280 35624 30308
rect 34011 30277 34023 30280
rect 33965 30271 34023 30277
rect 35618 30268 35624 30280
rect 35676 30268 35682 30320
rect 32125 30243 32183 30249
rect 32125 30209 32137 30243
rect 32171 30209 32183 30243
rect 32125 30203 32183 30209
rect 32401 30243 32459 30249
rect 32401 30209 32413 30243
rect 32447 30209 32459 30243
rect 32401 30203 32459 30209
rect 28316 30144 29868 30172
rect 28316 30132 28322 30144
rect 29914 30132 29920 30184
rect 29972 30172 29978 30184
rect 30009 30175 30067 30181
rect 30009 30172 30021 30175
rect 29972 30144 30021 30172
rect 29972 30132 29978 30144
rect 30009 30141 30021 30144
rect 30055 30141 30067 30175
rect 30282 30172 30288 30184
rect 30243 30144 30288 30172
rect 30009 30135 30067 30141
rect 30282 30132 30288 30144
rect 30340 30132 30346 30184
rect 30466 30132 30472 30184
rect 30524 30172 30530 30184
rect 31573 30175 31631 30181
rect 31573 30172 31585 30175
rect 30524 30144 31585 30172
rect 30524 30132 30530 30144
rect 31573 30141 31585 30144
rect 31619 30141 31631 30175
rect 32140 30172 32168 30203
rect 32490 30200 32496 30252
rect 32548 30240 32554 30252
rect 32861 30243 32919 30249
rect 32861 30240 32873 30243
rect 32548 30212 32873 30240
rect 32548 30200 32554 30212
rect 32861 30209 32873 30212
rect 32907 30209 32919 30243
rect 33042 30240 33048 30252
rect 33003 30212 33048 30240
rect 32861 30203 32919 30209
rect 33042 30200 33048 30212
rect 33100 30200 33106 30252
rect 34146 30240 34152 30252
rect 34107 30212 34152 30240
rect 34146 30200 34152 30212
rect 34204 30240 34210 30252
rect 34885 30243 34943 30249
rect 34885 30240 34897 30243
rect 34204 30212 34897 30240
rect 34204 30200 34210 30212
rect 34885 30209 34897 30212
rect 34931 30209 34943 30243
rect 36262 30240 36268 30252
rect 36223 30212 36268 30240
rect 34885 30203 34943 30209
rect 36262 30200 36268 30212
rect 36320 30200 36326 30252
rect 37461 30243 37519 30249
rect 37461 30209 37473 30243
rect 37507 30240 37519 30243
rect 37918 30240 37924 30252
rect 37507 30212 37924 30240
rect 37507 30209 37519 30212
rect 37461 30203 37519 30209
rect 37918 30200 37924 30212
rect 37976 30200 37982 30252
rect 34425 30175 34483 30181
rect 34425 30172 34437 30175
rect 32140 30144 34437 30172
rect 31573 30135 31631 30141
rect 34425 30141 34437 30144
rect 34471 30172 34483 30175
rect 35161 30175 35219 30181
rect 35161 30172 35173 30175
rect 34471 30144 35173 30172
rect 34471 30141 34483 30144
rect 34425 30135 34483 30141
rect 35161 30141 35173 30144
rect 35207 30141 35219 30175
rect 36170 30172 36176 30184
rect 36131 30144 36176 30172
rect 35161 30135 35219 30141
rect 36170 30132 36176 30144
rect 36228 30132 36234 30184
rect 37366 30172 37372 30184
rect 37327 30144 37372 30172
rect 37366 30132 37372 30144
rect 37424 30132 37430 30184
rect 25455 30076 26464 30104
rect 27433 30107 27491 30113
rect 25455 30073 25467 30076
rect 25409 30067 25467 30073
rect 27433 30073 27445 30107
rect 27479 30104 27491 30107
rect 34333 30107 34391 30113
rect 27479 30076 28304 30104
rect 27479 30073 27491 30076
rect 27433 30067 27491 30073
rect 16574 30036 16580 30048
rect 16040 30008 16580 30036
rect 16574 29996 16580 30008
rect 16632 29996 16638 30048
rect 17770 29996 17776 30048
rect 17828 30036 17834 30048
rect 22646 30036 22652 30048
rect 17828 30008 22652 30036
rect 17828 29996 17834 30008
rect 22646 29996 22652 30008
rect 22704 29996 22710 30048
rect 22830 30036 22836 30048
rect 22791 30008 22836 30036
rect 22830 29996 22836 30008
rect 22888 29996 22894 30048
rect 22922 29996 22928 30048
rect 22980 30036 22986 30048
rect 23017 30039 23075 30045
rect 23017 30036 23029 30039
rect 22980 30008 23029 30036
rect 22980 29996 22986 30008
rect 23017 30005 23029 30008
rect 23063 30005 23075 30039
rect 23017 29999 23075 30005
rect 24673 30039 24731 30045
rect 24673 30005 24685 30039
rect 24719 30036 24731 30039
rect 28074 30036 28080 30048
rect 24719 30008 28080 30036
rect 24719 30005 24731 30008
rect 24673 29999 24731 30005
rect 28074 29996 28080 30008
rect 28132 29996 28138 30048
rect 28276 30036 28304 30076
rect 28460 30076 34284 30104
rect 28460 30036 28488 30076
rect 28276 30008 28488 30036
rect 28626 29996 28632 30048
rect 28684 30036 28690 30048
rect 28905 30039 28963 30045
rect 28905 30036 28917 30039
rect 28684 30008 28917 30036
rect 28684 29996 28690 30008
rect 28905 30005 28917 30008
rect 28951 30036 28963 30039
rect 30926 30036 30932 30048
rect 28951 30008 30932 30036
rect 28951 30005 28963 30008
rect 28905 29999 28963 30005
rect 30926 29996 30932 30008
rect 30984 29996 30990 30048
rect 32125 30039 32183 30045
rect 32125 30005 32137 30039
rect 32171 30036 32183 30039
rect 32306 30036 32312 30048
rect 32171 30008 32312 30036
rect 32171 30005 32183 30008
rect 32125 29999 32183 30005
rect 32306 29996 32312 30008
rect 32364 29996 32370 30048
rect 32861 30039 32919 30045
rect 32861 30005 32873 30039
rect 32907 30036 32919 30039
rect 33962 30036 33968 30048
rect 32907 30008 33968 30036
rect 32907 30005 32919 30008
rect 32861 29999 32919 30005
rect 33962 29996 33968 30008
rect 34020 29996 34026 30048
rect 34256 30036 34284 30076
rect 34333 30073 34345 30107
rect 34379 30104 34391 30107
rect 34790 30104 34796 30116
rect 34379 30076 34796 30104
rect 34379 30073 34391 30076
rect 34333 30067 34391 30073
rect 34790 30064 34796 30076
rect 34848 30104 34854 30116
rect 34977 30107 35035 30113
rect 34977 30104 34989 30107
rect 34848 30076 34989 30104
rect 34848 30064 34854 30076
rect 34977 30073 34989 30076
rect 35023 30073 35035 30107
rect 37826 30104 37832 30116
rect 37787 30076 37832 30104
rect 34977 30067 35035 30073
rect 37826 30064 37832 30076
rect 37884 30064 37890 30116
rect 35894 30036 35900 30048
rect 34256 30008 35900 30036
rect 35894 29996 35900 30008
rect 35952 29996 35958 30048
rect 36538 30036 36544 30048
rect 36499 30008 36544 30036
rect 36538 29996 36544 30008
rect 36596 29996 36602 30048
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 15933 29835 15991 29841
rect 15933 29801 15945 29835
rect 15979 29832 15991 29835
rect 17034 29832 17040 29844
rect 15979 29804 17040 29832
rect 15979 29801 15991 29804
rect 15933 29795 15991 29801
rect 17034 29792 17040 29804
rect 17092 29792 17098 29844
rect 18046 29832 18052 29844
rect 18007 29804 18052 29832
rect 18046 29792 18052 29804
rect 18104 29792 18110 29844
rect 18325 29835 18383 29841
rect 18325 29801 18337 29835
rect 18371 29832 18383 29835
rect 19334 29832 19340 29844
rect 18371 29804 19340 29832
rect 18371 29801 18383 29804
rect 18325 29795 18383 29801
rect 19334 29792 19340 29804
rect 19392 29792 19398 29844
rect 19981 29835 20039 29841
rect 19981 29801 19993 29835
rect 20027 29832 20039 29835
rect 20070 29832 20076 29844
rect 20027 29804 20076 29832
rect 20027 29801 20039 29804
rect 19981 29795 20039 29801
rect 20070 29792 20076 29804
rect 20128 29792 20134 29844
rect 21266 29832 21272 29844
rect 21227 29804 21272 29832
rect 21266 29792 21272 29804
rect 21324 29832 21330 29844
rect 22830 29832 22836 29844
rect 21324 29804 22836 29832
rect 21324 29792 21330 29804
rect 22830 29792 22836 29804
rect 22888 29792 22894 29844
rect 22925 29835 22983 29841
rect 22925 29801 22937 29835
rect 22971 29832 22983 29835
rect 23014 29832 23020 29844
rect 22971 29804 23020 29832
rect 22971 29801 22983 29804
rect 22925 29795 22983 29801
rect 23014 29792 23020 29804
rect 23072 29792 23078 29844
rect 24581 29835 24639 29841
rect 24581 29801 24593 29835
rect 24627 29832 24639 29835
rect 24627 29804 24716 29832
rect 24627 29801 24639 29804
rect 24581 29795 24639 29801
rect 22462 29724 22468 29776
rect 22520 29764 22526 29776
rect 24688 29764 24716 29804
rect 25222 29792 25228 29844
rect 25280 29832 25286 29844
rect 26329 29835 26387 29841
rect 25280 29804 25820 29832
rect 25280 29792 25286 29804
rect 25038 29764 25044 29776
rect 22520 29736 24624 29764
rect 24688 29736 25044 29764
rect 22520 29724 22526 29736
rect 16022 29696 16028 29708
rect 15580 29668 16028 29696
rect 15580 29637 15608 29668
rect 16022 29656 16028 29668
rect 16080 29696 16086 29708
rect 16669 29699 16727 29705
rect 16669 29696 16681 29699
rect 16080 29668 16681 29696
rect 16080 29656 16086 29668
rect 16669 29665 16681 29668
rect 16715 29665 16727 29699
rect 16669 29659 16727 29665
rect 17402 29656 17408 29708
rect 17460 29696 17466 29708
rect 24210 29696 24216 29708
rect 17460 29668 24216 29696
rect 17460 29656 17466 29668
rect 15565 29631 15623 29637
rect 15565 29597 15577 29631
rect 15611 29597 15623 29631
rect 15565 29591 15623 29597
rect 16393 29631 16451 29637
rect 16393 29597 16405 29631
rect 16439 29628 16451 29631
rect 16574 29628 16580 29640
rect 16439 29600 16580 29628
rect 16439 29597 16451 29600
rect 16393 29591 16451 29597
rect 16574 29588 16580 29600
rect 16632 29588 16638 29640
rect 17954 29628 17960 29640
rect 17915 29600 17960 29628
rect 17954 29588 17960 29600
rect 18012 29588 18018 29640
rect 18141 29631 18199 29637
rect 18141 29597 18153 29631
rect 18187 29628 18199 29631
rect 18230 29628 18236 29640
rect 18187 29600 18236 29628
rect 18187 29597 18199 29600
rect 18141 29591 18199 29597
rect 18230 29588 18236 29600
rect 18288 29628 18294 29640
rect 21082 29628 21088 29640
rect 18288 29600 20392 29628
rect 21043 29600 21088 29628
rect 18288 29588 18294 29600
rect 15470 29520 15476 29572
rect 15528 29560 15534 29572
rect 15749 29563 15807 29569
rect 15749 29560 15761 29563
rect 15528 29532 15761 29560
rect 15528 29520 15534 29532
rect 15749 29529 15761 29532
rect 15795 29560 15807 29563
rect 15838 29560 15844 29572
rect 15795 29532 15844 29560
rect 15795 29529 15807 29532
rect 15749 29523 15807 29529
rect 15838 29520 15844 29532
rect 15896 29520 15902 29572
rect 16114 29520 16120 29572
rect 16172 29560 16178 29572
rect 19797 29563 19855 29569
rect 19797 29560 19809 29563
rect 16172 29532 19809 29560
rect 16172 29520 16178 29532
rect 19797 29529 19809 29532
rect 19843 29560 19855 29563
rect 20254 29560 20260 29572
rect 19843 29532 20260 29560
rect 19843 29529 19855 29532
rect 19797 29523 19855 29529
rect 20254 29520 20260 29532
rect 20312 29520 20318 29572
rect 20364 29560 20392 29600
rect 21082 29588 21088 29600
rect 21140 29588 21146 29640
rect 22649 29631 22707 29637
rect 22649 29628 22661 29631
rect 21192 29600 22661 29628
rect 21192 29560 21220 29600
rect 22649 29597 22661 29600
rect 22695 29628 22707 29631
rect 22738 29628 22744 29640
rect 22695 29600 22744 29628
rect 22695 29597 22707 29600
rect 22649 29591 22707 29597
rect 22738 29588 22744 29600
rect 22796 29588 22802 29640
rect 23382 29628 23388 29640
rect 23343 29600 23388 29628
rect 23382 29588 23388 29600
rect 23440 29588 23446 29640
rect 23584 29637 23612 29668
rect 24210 29656 24216 29668
rect 24268 29696 24274 29708
rect 24489 29699 24547 29705
rect 24489 29696 24501 29699
rect 24268 29668 24501 29696
rect 24268 29656 24274 29668
rect 24489 29665 24501 29668
rect 24535 29665 24547 29699
rect 24489 29659 24547 29665
rect 23569 29631 23627 29637
rect 23569 29597 23581 29631
rect 23615 29597 23627 29631
rect 23569 29591 23627 29597
rect 24397 29631 24455 29637
rect 24397 29597 24409 29631
rect 24443 29597 24455 29631
rect 24397 29591 24455 29597
rect 20364 29532 21220 29560
rect 22094 29520 22100 29572
rect 22152 29560 22158 29572
rect 22373 29563 22431 29569
rect 22373 29560 22385 29563
rect 22152 29532 22385 29560
rect 22152 29520 22158 29532
rect 22373 29529 22385 29532
rect 22419 29529 22431 29563
rect 22373 29523 22431 29529
rect 22557 29563 22615 29569
rect 22557 29529 22569 29563
rect 22603 29560 22615 29563
rect 23400 29560 23428 29588
rect 24118 29560 24124 29572
rect 22603 29532 23336 29560
rect 23400 29532 24124 29560
rect 22603 29529 22615 29532
rect 22557 29523 22615 29529
rect 19978 29452 19984 29504
rect 20036 29501 20042 29504
rect 20036 29495 20055 29501
rect 20043 29461 20055 29495
rect 20162 29492 20168 29504
rect 20123 29464 20168 29492
rect 20036 29455 20055 29461
rect 20036 29452 20042 29455
rect 20162 29452 20168 29464
rect 20220 29452 20226 29504
rect 22462 29452 22468 29504
rect 22520 29492 22526 29504
rect 22741 29495 22799 29501
rect 22741 29492 22753 29495
rect 22520 29464 22753 29492
rect 22520 29452 22526 29464
rect 22741 29461 22753 29464
rect 22787 29461 22799 29495
rect 23308 29492 23336 29532
rect 24118 29520 24124 29532
rect 24176 29560 24182 29572
rect 24412 29560 24440 29591
rect 24176 29532 24440 29560
rect 24596 29560 24624 29736
rect 25038 29724 25044 29736
rect 25096 29764 25102 29776
rect 25682 29764 25688 29776
rect 25096 29736 25544 29764
rect 25643 29736 25688 29764
rect 25096 29724 25102 29736
rect 24670 29656 24676 29708
rect 24728 29696 24734 29708
rect 25222 29696 25228 29708
rect 24728 29668 24773 29696
rect 25148 29668 25228 29696
rect 24728 29656 24734 29668
rect 24762 29588 24768 29640
rect 24820 29628 24826 29640
rect 25148 29628 25176 29668
rect 25222 29656 25228 29668
rect 25280 29656 25286 29708
rect 25406 29696 25412 29708
rect 25367 29668 25412 29696
rect 25406 29656 25412 29668
rect 25464 29656 25470 29708
rect 25516 29696 25544 29736
rect 25682 29724 25688 29736
rect 25740 29724 25746 29776
rect 25792 29764 25820 29804
rect 26329 29801 26341 29835
rect 26375 29832 26387 29835
rect 28994 29832 29000 29844
rect 26375 29804 26648 29832
rect 26375 29801 26387 29804
rect 26329 29795 26387 29801
rect 26513 29767 26571 29773
rect 26513 29764 26525 29767
rect 25792 29736 26525 29764
rect 26513 29733 26525 29736
rect 26559 29733 26571 29767
rect 26513 29727 26571 29733
rect 26620 29696 26648 29804
rect 28966 29792 29000 29832
rect 29052 29832 29058 29844
rect 29362 29832 29368 29844
rect 29052 29804 29368 29832
rect 29052 29792 29058 29804
rect 29362 29792 29368 29804
rect 29420 29832 29426 29844
rect 34698 29832 34704 29844
rect 29420 29804 34704 29832
rect 29420 29792 29426 29804
rect 34698 29792 34704 29804
rect 34756 29792 34762 29844
rect 36081 29835 36139 29841
rect 36081 29801 36093 29835
rect 36127 29832 36139 29835
rect 37366 29832 37372 29844
rect 36127 29804 37372 29832
rect 36127 29801 36139 29804
rect 36081 29795 36139 29801
rect 37366 29792 37372 29804
rect 37424 29792 37430 29844
rect 28966 29764 28994 29792
rect 33594 29764 33600 29776
rect 25516 29668 26648 29696
rect 27632 29736 28994 29764
rect 29748 29736 33600 29764
rect 25314 29628 25320 29640
rect 24820 29600 25176 29628
rect 25275 29600 25320 29628
rect 24820 29588 24826 29600
rect 25314 29588 25320 29600
rect 25372 29588 25378 29640
rect 27632 29628 27660 29736
rect 27801 29699 27859 29705
rect 27801 29665 27813 29699
rect 27847 29696 27859 29699
rect 28902 29696 28908 29708
rect 27847 29668 28908 29696
rect 27847 29665 27859 29668
rect 27801 29659 27859 29665
rect 28902 29656 28908 29668
rect 28960 29656 28966 29708
rect 29086 29656 29092 29708
rect 29144 29696 29150 29708
rect 29748 29696 29776 29736
rect 33594 29724 33600 29736
rect 33652 29724 33658 29776
rect 33689 29767 33747 29773
rect 33689 29733 33701 29767
rect 33735 29764 33747 29767
rect 34146 29764 34152 29776
rect 33735 29736 34152 29764
rect 33735 29733 33747 29736
rect 33689 29727 33747 29733
rect 34146 29724 34152 29736
rect 34204 29724 34210 29776
rect 36262 29764 36268 29776
rect 34716 29736 36268 29764
rect 29144 29668 29776 29696
rect 30193 29699 30251 29705
rect 29144 29656 29150 29668
rect 30193 29665 30205 29699
rect 30239 29696 30251 29699
rect 30650 29696 30656 29708
rect 30239 29668 30656 29696
rect 30239 29665 30251 29668
rect 30193 29659 30251 29665
rect 30650 29656 30656 29668
rect 30708 29696 30714 29708
rect 31846 29696 31852 29708
rect 30708 29668 31754 29696
rect 31807 29668 31852 29696
rect 30708 29656 30714 29668
rect 26068 29600 27660 29628
rect 26068 29560 26096 29600
rect 28074 29588 28080 29640
rect 28132 29588 28138 29640
rect 28629 29631 28687 29637
rect 28629 29597 28641 29631
rect 28675 29628 28687 29631
rect 31021 29631 31079 29637
rect 28675 29600 30972 29628
rect 28675 29597 28687 29600
rect 28629 29591 28687 29597
rect 24596 29532 26096 29560
rect 24176 29520 24182 29532
rect 26142 29520 26148 29572
rect 26200 29560 26206 29572
rect 29178 29560 29184 29572
rect 26200 29532 29184 29560
rect 26200 29520 26206 29532
rect 29178 29520 29184 29532
rect 29236 29520 29242 29572
rect 30006 29560 30012 29572
rect 29967 29532 30012 29560
rect 30006 29520 30012 29532
rect 30064 29520 30070 29572
rect 30837 29563 30895 29569
rect 30837 29529 30849 29563
rect 30883 29529 30895 29563
rect 30944 29560 30972 29600
rect 31021 29597 31033 29631
rect 31067 29628 31079 29631
rect 31202 29628 31208 29640
rect 31067 29600 31208 29628
rect 31067 29597 31079 29600
rect 31021 29591 31079 29597
rect 31202 29588 31208 29600
rect 31260 29588 31266 29640
rect 31726 29628 31754 29668
rect 31846 29656 31852 29668
rect 31904 29656 31910 29708
rect 32125 29699 32183 29705
rect 32125 29665 32137 29699
rect 32171 29696 32183 29699
rect 32214 29696 32220 29708
rect 32171 29668 32220 29696
rect 32171 29665 32183 29668
rect 32125 29659 32183 29665
rect 32214 29656 32220 29668
rect 32272 29656 32278 29708
rect 32858 29696 32864 29708
rect 32416 29668 32864 29696
rect 32416 29628 32444 29668
rect 32858 29656 32864 29668
rect 32916 29656 32922 29708
rect 33226 29696 33232 29708
rect 33187 29668 33232 29696
rect 33226 29656 33232 29668
rect 33284 29656 33290 29708
rect 34716 29696 34744 29736
rect 36262 29724 36268 29736
rect 36320 29724 36326 29776
rect 33704 29668 34744 29696
rect 31726 29600 32444 29628
rect 32490 29588 32496 29640
rect 32548 29628 32554 29640
rect 33321 29631 33379 29637
rect 33321 29628 33333 29631
rect 32548 29600 33333 29628
rect 32548 29588 32554 29600
rect 33321 29597 33333 29600
rect 33367 29597 33379 29631
rect 33321 29591 33379 29597
rect 33704 29560 33732 29668
rect 34790 29656 34796 29708
rect 34848 29696 34854 29708
rect 34848 29668 35572 29696
rect 34848 29656 34854 29668
rect 33962 29588 33968 29640
rect 34020 29628 34026 29640
rect 34514 29628 34520 29640
rect 34020 29600 34520 29628
rect 34020 29588 34026 29600
rect 34514 29588 34520 29600
rect 34572 29588 34578 29640
rect 34698 29628 34704 29640
rect 34659 29600 34704 29628
rect 34698 29588 34704 29600
rect 34756 29588 34762 29640
rect 34885 29631 34943 29637
rect 34885 29597 34897 29631
rect 34931 29628 34943 29631
rect 34974 29628 34980 29640
rect 34931 29600 34980 29628
rect 34931 29597 34943 29600
rect 34885 29591 34943 29597
rect 34974 29588 34980 29600
rect 35032 29588 35038 29640
rect 35544 29637 35572 29668
rect 35345 29631 35403 29637
rect 35345 29597 35357 29631
rect 35391 29597 35403 29631
rect 35345 29591 35403 29597
rect 35529 29631 35587 29637
rect 35529 29597 35541 29631
rect 35575 29597 35587 29631
rect 35529 29591 35587 29597
rect 30944 29532 33732 29560
rect 30837 29523 30895 29529
rect 23474 29492 23480 29504
rect 23308 29464 23480 29492
rect 22741 29455 22799 29461
rect 23474 29452 23480 29464
rect 23532 29452 23538 29504
rect 23661 29495 23719 29501
rect 23661 29461 23673 29495
rect 23707 29492 23719 29495
rect 23750 29492 23756 29504
rect 23707 29464 23756 29492
rect 23707 29461 23719 29464
rect 23661 29455 23719 29461
rect 23750 29452 23756 29464
rect 23808 29492 23814 29504
rect 24026 29492 24032 29504
rect 23808 29464 24032 29492
rect 23808 29452 23814 29464
rect 24026 29452 24032 29464
rect 24084 29452 24090 29504
rect 24578 29452 24584 29504
rect 24636 29492 24642 29504
rect 26345 29495 26403 29501
rect 26345 29492 26357 29495
rect 24636 29464 26357 29492
rect 24636 29452 24642 29464
rect 26345 29461 26357 29464
rect 26391 29461 26403 29495
rect 26345 29455 26403 29461
rect 27246 29452 27252 29504
rect 27304 29492 27310 29504
rect 28166 29492 28172 29504
rect 27304 29464 28172 29492
rect 27304 29452 27310 29464
rect 28166 29452 28172 29464
rect 28224 29452 28230 29504
rect 29270 29452 29276 29504
rect 29328 29492 29334 29504
rect 29914 29492 29920 29504
rect 29328 29464 29920 29492
rect 29328 29452 29334 29464
rect 29914 29452 29920 29464
rect 29972 29492 29978 29504
rect 30098 29492 30104 29504
rect 29972 29464 30104 29492
rect 29972 29452 29978 29464
rect 30098 29452 30104 29464
rect 30156 29452 30162 29504
rect 30852 29492 30880 29523
rect 33778 29520 33784 29572
rect 33836 29560 33842 29572
rect 35360 29560 35388 29591
rect 35618 29588 35624 29640
rect 35676 29628 35682 29640
rect 36081 29631 36139 29637
rect 36081 29628 36093 29631
rect 35676 29600 36093 29628
rect 35676 29588 35682 29600
rect 36081 29597 36093 29600
rect 36127 29597 36139 29631
rect 36081 29591 36139 29597
rect 36170 29588 36176 29640
rect 36228 29628 36234 29640
rect 36357 29631 36415 29637
rect 36357 29628 36369 29631
rect 36228 29600 36369 29628
rect 36228 29588 36234 29600
rect 36357 29597 36369 29600
rect 36403 29597 36415 29631
rect 36357 29591 36415 29597
rect 36262 29560 36268 29572
rect 33836 29532 35388 29560
rect 36223 29532 36268 29560
rect 33836 29520 33842 29532
rect 36262 29520 36268 29532
rect 36320 29520 36326 29572
rect 32214 29492 32220 29504
rect 30852 29464 32220 29492
rect 32214 29452 32220 29464
rect 32272 29452 32278 29504
rect 32950 29452 32956 29504
rect 33008 29492 33014 29504
rect 34793 29495 34851 29501
rect 34793 29492 34805 29495
rect 33008 29464 34805 29492
rect 33008 29452 33014 29464
rect 34793 29461 34805 29464
rect 34839 29461 34851 29495
rect 34793 29455 34851 29461
rect 34882 29452 34888 29504
rect 34940 29492 34946 29504
rect 35437 29495 35495 29501
rect 35437 29492 35449 29495
rect 34940 29464 35449 29492
rect 34940 29452 34946 29464
rect 35437 29461 35449 29464
rect 35483 29461 35495 29495
rect 35437 29455 35495 29461
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 17402 29288 17408 29300
rect 17363 29260 17408 29288
rect 17402 29248 17408 29260
rect 17460 29248 17466 29300
rect 17770 29288 17776 29300
rect 17731 29260 17776 29288
rect 17770 29248 17776 29260
rect 17828 29248 17834 29300
rect 18248 29260 20116 29288
rect 15838 29180 15844 29232
rect 15896 29220 15902 29232
rect 16761 29223 16819 29229
rect 16761 29220 16773 29223
rect 15896 29192 16773 29220
rect 15896 29180 15902 29192
rect 16761 29189 16773 29192
rect 16807 29189 16819 29223
rect 16942 29220 16948 29232
rect 16903 29192 16948 29220
rect 16761 29183 16819 29189
rect 16942 29180 16948 29192
rect 17000 29180 17006 29232
rect 15933 29155 15991 29161
rect 15933 29121 15945 29155
rect 15979 29121 15991 29155
rect 16114 29152 16120 29164
rect 16075 29124 16120 29152
rect 15933 29115 15991 29121
rect 15948 29084 15976 29115
rect 16114 29112 16120 29124
rect 16172 29112 16178 29164
rect 17586 29152 17592 29164
rect 17547 29124 17592 29152
rect 17586 29112 17592 29124
rect 17644 29112 17650 29164
rect 17862 29152 17868 29164
rect 17823 29124 17868 29152
rect 17862 29112 17868 29124
rect 17920 29112 17926 29164
rect 18248 29096 18276 29260
rect 19978 29220 19984 29232
rect 19720 29192 19984 29220
rect 19720 29164 19748 29192
rect 19978 29180 19984 29192
rect 20036 29180 20042 29232
rect 20088 29164 20116 29260
rect 22186 29248 22192 29300
rect 22244 29288 22250 29300
rect 23017 29291 23075 29297
rect 23017 29288 23029 29291
rect 22244 29260 23029 29288
rect 22244 29248 22250 29260
rect 23017 29257 23029 29260
rect 23063 29257 23075 29291
rect 24762 29288 24768 29300
rect 23017 29251 23075 29257
rect 23952 29260 24768 29288
rect 21082 29180 21088 29232
rect 21140 29220 21146 29232
rect 21140 29192 23152 29220
rect 21140 29180 21146 29192
rect 18325 29155 18383 29161
rect 18325 29121 18337 29155
rect 18371 29121 18383 29155
rect 18506 29152 18512 29164
rect 18467 29124 18512 29152
rect 18325 29115 18383 29121
rect 18230 29084 18236 29096
rect 15948 29056 18236 29084
rect 18230 29044 18236 29056
rect 18288 29044 18294 29096
rect 18340 29084 18368 29115
rect 18506 29112 18512 29124
rect 18564 29112 18570 29164
rect 19521 29155 19579 29161
rect 19521 29121 19533 29155
rect 19567 29121 19579 29155
rect 19702 29152 19708 29164
rect 19663 29124 19708 29152
rect 19521 29115 19579 29121
rect 18598 29084 18604 29096
rect 18340 29056 18604 29084
rect 18598 29044 18604 29056
rect 18656 29044 18662 29096
rect 19536 29084 19564 29115
rect 19702 29112 19708 29124
rect 19760 29112 19766 29164
rect 19889 29155 19947 29161
rect 19889 29121 19901 29155
rect 19935 29152 19947 29155
rect 20070 29152 20076 29164
rect 19935 29124 20076 29152
rect 19935 29121 19947 29124
rect 19889 29115 19947 29121
rect 20070 29112 20076 29124
rect 20128 29112 20134 29164
rect 20254 29152 20260 29164
rect 20215 29124 20260 29152
rect 20254 29112 20260 29124
rect 20312 29112 20318 29164
rect 20346 29112 20352 29164
rect 20404 29152 20410 29164
rect 20717 29155 20775 29161
rect 20717 29152 20729 29155
rect 20404 29124 20729 29152
rect 20404 29112 20410 29124
rect 20717 29121 20729 29124
rect 20763 29121 20775 29155
rect 20717 29115 20775 29121
rect 20898 29112 20904 29164
rect 20956 29152 20962 29164
rect 21910 29152 21916 29164
rect 20956 29124 21916 29152
rect 20956 29112 20962 29124
rect 21910 29112 21916 29124
rect 21968 29152 21974 29164
rect 22281 29155 22339 29161
rect 22281 29152 22293 29155
rect 21968 29124 22293 29152
rect 21968 29112 21974 29124
rect 22281 29121 22293 29124
rect 22327 29121 22339 29155
rect 22281 29115 22339 29121
rect 22925 29155 22983 29161
rect 22925 29121 22937 29155
rect 22971 29152 22983 29155
rect 23014 29152 23020 29164
rect 22971 29124 23020 29152
rect 22971 29121 22983 29124
rect 22925 29115 22983 29121
rect 23014 29112 23020 29124
rect 23072 29112 23078 29164
rect 23124 29161 23152 29192
rect 23109 29155 23167 29161
rect 23109 29121 23121 29155
rect 23155 29121 23167 29155
rect 23842 29152 23848 29164
rect 23803 29124 23848 29152
rect 23109 29115 23167 29121
rect 23842 29112 23848 29124
rect 23900 29112 23906 29164
rect 23952 29161 23980 29260
rect 24762 29248 24768 29260
rect 24820 29248 24826 29300
rect 26142 29288 26148 29300
rect 24872 29260 26148 29288
rect 24103 29161 24109 29164
rect 23937 29155 23995 29161
rect 23937 29121 23949 29155
rect 23983 29121 23995 29155
rect 23937 29115 23995 29121
rect 24080 29155 24109 29161
rect 24080 29121 24092 29155
rect 24080 29115 24109 29121
rect 24103 29112 24109 29115
rect 24161 29112 24167 29164
rect 24210 29112 24216 29164
rect 24268 29161 24274 29164
rect 24872 29161 24900 29260
rect 26142 29248 26148 29260
rect 26200 29248 26206 29300
rect 27433 29291 27491 29297
rect 27433 29257 27445 29291
rect 27479 29288 27491 29291
rect 27614 29288 27620 29300
rect 27479 29260 27620 29288
rect 27479 29257 27491 29260
rect 27433 29251 27491 29257
rect 27614 29248 27620 29260
rect 27672 29248 27678 29300
rect 28074 29288 28080 29300
rect 28035 29260 28080 29288
rect 28074 29248 28080 29260
rect 28132 29248 28138 29300
rect 28718 29288 28724 29300
rect 28776 29297 28782 29300
rect 28776 29291 28795 29297
rect 28184 29260 28724 29288
rect 25222 29180 25228 29232
rect 25280 29220 25286 29232
rect 25280 29192 27108 29220
rect 25280 29180 25286 29192
rect 24268 29155 24281 29161
rect 24269 29152 24281 29155
rect 24857 29155 24915 29161
rect 24857 29152 24869 29155
rect 24269 29124 24313 29152
rect 24504 29124 24869 29152
rect 24269 29121 24281 29124
rect 24268 29115 24281 29121
rect 24268 29112 24274 29115
rect 21726 29084 21732 29096
rect 19536 29056 21732 29084
rect 21726 29044 21732 29056
rect 21784 29044 21790 29096
rect 24504 29084 24532 29124
rect 24857 29121 24869 29124
rect 24903 29121 24915 29155
rect 25038 29152 25044 29164
rect 24999 29124 25044 29152
rect 24857 29115 24915 29121
rect 25038 29112 25044 29124
rect 25096 29112 25102 29164
rect 25133 29155 25191 29161
rect 25133 29121 25145 29155
rect 25179 29121 25191 29155
rect 25133 29115 25191 29121
rect 26053 29155 26111 29161
rect 26053 29121 26065 29155
rect 26099 29152 26111 29155
rect 26510 29152 26516 29164
rect 26099 29124 26516 29152
rect 26099 29121 26111 29124
rect 26053 29115 26111 29121
rect 22480 29056 24532 29084
rect 16025 29019 16083 29025
rect 16025 28985 16037 29019
rect 16071 29016 16083 29019
rect 20714 29016 20720 29028
rect 16071 28988 20720 29016
rect 16071 28985 16083 28988
rect 16025 28979 16083 28985
rect 20714 28976 20720 28988
rect 20772 28976 20778 29028
rect 22480 29025 22508 29056
rect 24578 29044 24584 29096
rect 24636 29084 24642 29096
rect 25148 29084 25176 29115
rect 24636 29056 25176 29084
rect 24636 29044 24642 29056
rect 22465 29019 22523 29025
rect 22465 28985 22477 29019
rect 22511 28985 22523 29019
rect 22465 28979 22523 28985
rect 24394 28976 24400 29028
rect 24452 29016 24458 29028
rect 26068 29016 26096 29115
rect 26510 29112 26516 29124
rect 26568 29152 26574 29164
rect 27080 29152 27108 29192
rect 27154 29180 27160 29232
rect 27212 29220 27218 29232
rect 28184 29220 28212 29260
rect 28718 29248 28724 29260
rect 28783 29257 28795 29291
rect 30006 29288 30012 29300
rect 28776 29251 28795 29257
rect 28828 29260 30012 29288
rect 28776 29248 28782 29251
rect 28534 29220 28540 29232
rect 27212 29192 28212 29220
rect 28447 29192 28540 29220
rect 27212 29180 27218 29192
rect 28534 29180 28540 29192
rect 28592 29220 28598 29232
rect 28828 29220 28856 29260
rect 30006 29248 30012 29260
rect 30064 29248 30070 29300
rect 31297 29291 31355 29297
rect 31297 29257 31309 29291
rect 31343 29288 31355 29291
rect 31938 29288 31944 29300
rect 31343 29260 31944 29288
rect 31343 29257 31355 29260
rect 31297 29251 31355 29257
rect 31938 29248 31944 29260
rect 31996 29248 32002 29300
rect 32306 29248 32312 29300
rect 32364 29297 32370 29300
rect 32364 29291 32383 29297
rect 32371 29257 32383 29291
rect 32364 29251 32383 29257
rect 32493 29291 32551 29297
rect 32493 29257 32505 29291
rect 32539 29257 32551 29291
rect 32493 29251 32551 29257
rect 32364 29248 32370 29251
rect 28592 29192 28856 29220
rect 28592 29180 28598 29192
rect 28902 29180 28908 29232
rect 28960 29220 28966 29232
rect 29086 29220 29092 29232
rect 28960 29192 29092 29220
rect 28960 29180 28966 29192
rect 29086 29180 29092 29192
rect 29144 29180 29150 29232
rect 29641 29223 29699 29229
rect 29641 29220 29653 29223
rect 29564 29192 29653 29220
rect 29270 29152 29276 29164
rect 26568 29124 27016 29152
rect 27080 29124 29276 29152
rect 26568 29112 26574 29124
rect 26237 29087 26295 29093
rect 26237 29053 26249 29087
rect 26283 29084 26295 29087
rect 26602 29084 26608 29096
rect 26283 29056 26608 29084
rect 26283 29053 26295 29056
rect 26237 29047 26295 29053
rect 26602 29044 26608 29056
rect 26660 29044 26666 29096
rect 24452 28988 26096 29016
rect 26988 29016 27016 29124
rect 29270 29112 29276 29124
rect 29328 29112 29334 29164
rect 29454 29152 29460 29164
rect 29415 29124 29460 29152
rect 29454 29112 29460 29124
rect 29512 29112 29518 29164
rect 27246 29044 27252 29096
rect 27304 29084 27310 29096
rect 27801 29087 27859 29093
rect 27801 29084 27813 29087
rect 27304 29056 27813 29084
rect 27304 29044 27310 29056
rect 27801 29053 27813 29056
rect 27847 29053 27859 29087
rect 27801 29047 27859 29053
rect 27893 29087 27951 29093
rect 27893 29053 27905 29087
rect 27939 29053 27951 29087
rect 27893 29047 27951 29053
rect 27706 29016 27712 29028
rect 26988 28988 27712 29016
rect 24452 28976 24458 28988
rect 27706 28976 27712 28988
rect 27764 28976 27770 29028
rect 27908 29016 27936 29047
rect 29362 29044 29368 29096
rect 29420 29084 29426 29096
rect 29564 29084 29592 29192
rect 29641 29189 29653 29192
rect 29687 29189 29699 29223
rect 29641 29183 29699 29189
rect 32030 29180 32036 29232
rect 32088 29220 32094 29232
rect 32125 29223 32183 29229
rect 32125 29220 32137 29223
rect 32088 29192 32137 29220
rect 32088 29180 32094 29192
rect 32125 29189 32137 29192
rect 32171 29189 32183 29223
rect 32508 29220 32536 29251
rect 32674 29248 32680 29300
rect 32732 29288 32738 29300
rect 33042 29288 33048 29300
rect 32732 29260 33048 29288
rect 32732 29248 32738 29260
rect 33042 29248 33048 29260
rect 33100 29248 33106 29300
rect 33226 29288 33232 29300
rect 33187 29260 33232 29288
rect 33226 29248 33232 29260
rect 33284 29248 33290 29300
rect 34330 29248 34336 29300
rect 34388 29288 34394 29300
rect 34974 29288 34980 29300
rect 34388 29260 34980 29288
rect 34388 29248 34394 29260
rect 34974 29248 34980 29260
rect 35032 29248 35038 29300
rect 37918 29288 37924 29300
rect 37879 29260 37924 29288
rect 37918 29248 37924 29260
rect 37976 29248 37982 29300
rect 34790 29220 34796 29232
rect 32508 29192 34796 29220
rect 32125 29183 32183 29189
rect 34790 29180 34796 29192
rect 34848 29180 34854 29232
rect 36449 29223 36507 29229
rect 36449 29189 36461 29223
rect 36495 29220 36507 29223
rect 36538 29220 36544 29232
rect 36495 29192 36544 29220
rect 36495 29189 36507 29192
rect 36449 29183 36507 29189
rect 36538 29180 36544 29192
rect 36596 29180 36602 29232
rect 29733 29155 29791 29161
rect 29733 29121 29745 29155
rect 29779 29121 29791 29155
rect 29733 29115 29791 29121
rect 29825 29155 29883 29161
rect 29825 29121 29837 29155
rect 29871 29121 29883 29155
rect 29825 29115 29883 29121
rect 29420 29056 29592 29084
rect 29420 29044 29426 29056
rect 29638 29044 29644 29096
rect 29696 29084 29702 29096
rect 29748 29084 29776 29115
rect 29696 29056 29776 29084
rect 29840 29084 29868 29115
rect 30374 29112 30380 29164
rect 30432 29152 30438 29164
rect 30469 29155 30527 29161
rect 30469 29152 30481 29155
rect 30432 29124 30481 29152
rect 30432 29112 30438 29124
rect 30469 29121 30481 29124
rect 30515 29121 30527 29155
rect 30650 29152 30656 29164
rect 30611 29124 30656 29152
rect 30469 29115 30527 29121
rect 30650 29112 30656 29124
rect 30708 29112 30714 29164
rect 31202 29152 31208 29164
rect 31163 29124 31208 29152
rect 31202 29112 31208 29124
rect 31260 29112 31266 29164
rect 32950 29152 32956 29164
rect 32911 29124 32956 29152
rect 32950 29112 32956 29124
rect 33008 29112 33014 29164
rect 33870 29152 33876 29164
rect 33831 29124 33876 29152
rect 33870 29112 33876 29124
rect 33928 29112 33934 29164
rect 34698 29152 34704 29164
rect 34611 29124 34704 29152
rect 34698 29112 34704 29124
rect 34756 29152 34762 29164
rect 34882 29152 34888 29164
rect 34756 29124 34888 29152
rect 34756 29112 34762 29124
rect 34882 29112 34888 29124
rect 34940 29112 34946 29164
rect 35713 29155 35771 29161
rect 35713 29152 35725 29155
rect 35084 29124 35725 29152
rect 30098 29084 30104 29096
rect 29840 29056 30104 29084
rect 29696 29044 29702 29056
rect 30098 29044 30104 29056
rect 30156 29044 30162 29096
rect 33226 29084 33232 29096
rect 33187 29056 33232 29084
rect 33226 29044 33232 29056
rect 33284 29044 33290 29096
rect 33962 29084 33968 29096
rect 33923 29056 33968 29084
rect 33962 29044 33968 29056
rect 34020 29044 34026 29096
rect 34514 29044 34520 29096
rect 34572 29084 34578 29096
rect 34793 29087 34851 29093
rect 34793 29084 34805 29087
rect 34572 29056 34805 29084
rect 34572 29044 34578 29056
rect 34793 29053 34805 29056
rect 34839 29053 34851 29087
rect 34793 29047 34851 29053
rect 28442 29016 28448 29028
rect 27908 28988 28448 29016
rect 28442 28976 28448 28988
rect 28500 29016 28506 29028
rect 28905 29019 28963 29025
rect 28905 29016 28917 29019
rect 28500 28988 28917 29016
rect 28500 28976 28506 28988
rect 28905 28985 28917 28988
rect 28951 28985 28963 29019
rect 30558 29016 30564 29028
rect 28905 28979 28963 28985
rect 29932 28988 30236 29016
rect 30471 28988 30564 29016
rect 18414 28948 18420 28960
rect 18375 28920 18420 28948
rect 18414 28908 18420 28920
rect 18472 28908 18478 28960
rect 19242 28908 19248 28960
rect 19300 28948 19306 28960
rect 19521 28951 19579 28957
rect 19521 28948 19533 28951
rect 19300 28920 19533 28948
rect 19300 28908 19306 28920
rect 19521 28917 19533 28920
rect 19567 28917 19579 28951
rect 19521 28911 19579 28917
rect 20254 28908 20260 28960
rect 20312 28948 20318 28960
rect 20530 28948 20536 28960
rect 20312 28920 20536 28948
rect 20312 28908 20318 28920
rect 20530 28908 20536 28920
rect 20588 28908 20594 28960
rect 20809 28951 20867 28957
rect 20809 28917 20821 28951
rect 20855 28948 20867 28951
rect 20898 28948 20904 28960
rect 20855 28920 20904 28948
rect 20855 28917 20867 28920
rect 20809 28911 20867 28917
rect 20898 28908 20904 28920
rect 20956 28908 20962 28960
rect 23661 28951 23719 28957
rect 23661 28917 23673 28951
rect 23707 28948 23719 28951
rect 24578 28948 24584 28960
rect 23707 28920 24584 28948
rect 23707 28917 23719 28920
rect 23661 28911 23719 28917
rect 24578 28908 24584 28920
rect 24636 28908 24642 28960
rect 24673 28951 24731 28957
rect 24673 28917 24685 28951
rect 24719 28948 24731 28951
rect 24946 28948 24952 28960
rect 24719 28920 24952 28948
rect 24719 28917 24731 28920
rect 24673 28911 24731 28917
rect 24946 28908 24952 28920
rect 25004 28908 25010 28960
rect 25866 28908 25872 28960
rect 25924 28948 25930 28960
rect 28721 28951 28779 28957
rect 28721 28948 28733 28951
rect 25924 28920 28733 28948
rect 25924 28908 25930 28920
rect 28721 28917 28733 28920
rect 28767 28948 28779 28951
rect 29454 28948 29460 28960
rect 28767 28920 29460 28948
rect 28767 28917 28779 28920
rect 28721 28911 28779 28917
rect 29454 28908 29460 28920
rect 29512 28908 29518 28960
rect 29730 28908 29736 28960
rect 29788 28948 29794 28960
rect 29932 28948 29960 28988
rect 29788 28920 29960 28948
rect 30009 28951 30067 28957
rect 29788 28908 29794 28920
rect 30009 28917 30021 28951
rect 30055 28948 30067 28951
rect 30098 28948 30104 28960
rect 30055 28920 30104 28948
rect 30055 28917 30067 28920
rect 30009 28911 30067 28917
rect 30098 28908 30104 28920
rect 30156 28908 30162 28960
rect 30208 28948 30236 28988
rect 30558 28976 30564 28988
rect 30616 29016 30622 29028
rect 31202 29016 31208 29028
rect 30616 28988 31208 29016
rect 30616 28976 30622 28988
rect 31202 28976 31208 28988
rect 31260 28976 31266 29028
rect 32674 29016 32680 29028
rect 31726 28988 32680 29016
rect 31726 28948 31754 28988
rect 32674 28976 32680 28988
rect 32732 28976 32738 29028
rect 34146 28976 34152 29028
rect 34204 28976 34210 29028
rect 34241 29019 34299 29025
rect 34241 28985 34253 29019
rect 34287 29016 34299 29019
rect 34606 29016 34612 29028
rect 34287 28988 34612 29016
rect 34287 28985 34299 28988
rect 34241 28979 34299 28985
rect 34606 28976 34612 28988
rect 34664 28976 34670 29028
rect 35084 29025 35112 29124
rect 35713 29121 35725 29124
rect 35759 29121 35771 29155
rect 36630 29152 36636 29164
rect 36591 29124 36636 29152
rect 35713 29115 35771 29121
rect 36630 29112 36636 29124
rect 36688 29112 36694 29164
rect 36725 29155 36783 29161
rect 36725 29121 36737 29155
rect 36771 29121 36783 29155
rect 36725 29115 36783 29121
rect 35526 29084 35532 29096
rect 35487 29056 35532 29084
rect 35526 29044 35532 29056
rect 35584 29084 35590 29096
rect 36740 29084 36768 29115
rect 37274 29084 37280 29096
rect 35584 29056 36768 29084
rect 37235 29056 37280 29084
rect 35584 29044 35590 29056
rect 37274 29044 37280 29056
rect 37332 29044 37338 29096
rect 37458 29044 37464 29096
rect 37516 29084 37522 29096
rect 37645 29087 37703 29093
rect 37645 29084 37657 29087
rect 37516 29056 37657 29084
rect 37516 29044 37522 29056
rect 37645 29053 37657 29056
rect 37691 29053 37703 29087
rect 37645 29047 37703 29053
rect 37737 29087 37795 29093
rect 37737 29053 37749 29087
rect 37783 29053 37795 29087
rect 37737 29047 37795 29053
rect 35069 29019 35127 29025
rect 35069 28985 35081 29019
rect 35115 28985 35127 29019
rect 35069 28979 35127 28985
rect 36725 29019 36783 29025
rect 36725 28985 36737 29019
rect 36771 29016 36783 29019
rect 37752 29016 37780 29047
rect 37918 29016 37924 29028
rect 36771 28988 37924 29016
rect 36771 28985 36783 28988
rect 36725 28979 36783 28985
rect 37918 28976 37924 28988
rect 37976 28976 37982 29028
rect 30208 28920 31754 28948
rect 31846 28908 31852 28960
rect 31904 28948 31910 28960
rect 32309 28951 32367 28957
rect 32309 28948 32321 28951
rect 31904 28920 32321 28948
rect 31904 28908 31910 28920
rect 32309 28917 32321 28920
rect 32355 28917 32367 28951
rect 33042 28948 33048 28960
rect 33003 28920 33048 28948
rect 32309 28911 32367 28917
rect 33042 28908 33048 28920
rect 33100 28908 33106 28960
rect 34164 28948 34192 28976
rect 34422 28948 34428 28960
rect 34164 28920 34428 28948
rect 34422 28908 34428 28920
rect 34480 28908 34486 28960
rect 34790 28948 34796 28960
rect 34751 28920 34796 28948
rect 34790 28908 34796 28920
rect 34848 28908 34854 28960
rect 35894 28948 35900 28960
rect 35855 28920 35900 28948
rect 35894 28908 35900 28920
rect 35952 28908 35958 28960
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 15470 28744 15476 28756
rect 15431 28716 15476 28744
rect 15470 28704 15476 28716
rect 15528 28704 15534 28756
rect 16574 28704 16580 28756
rect 16632 28744 16638 28756
rect 16945 28747 17003 28753
rect 16945 28744 16957 28747
rect 16632 28716 16957 28744
rect 16632 28704 16638 28716
rect 16945 28713 16957 28716
rect 16991 28713 17003 28747
rect 16945 28707 17003 28713
rect 17218 28704 17224 28756
rect 17276 28744 17282 28756
rect 18509 28747 18567 28753
rect 18509 28744 18521 28747
rect 17276 28716 18521 28744
rect 17276 28704 17282 28716
rect 18509 28713 18521 28716
rect 18555 28744 18567 28747
rect 18555 28716 18828 28744
rect 18555 28713 18567 28716
rect 18509 28707 18567 28713
rect 18693 28679 18751 28685
rect 18693 28645 18705 28679
rect 18739 28645 18751 28679
rect 18800 28676 18828 28716
rect 19150 28704 19156 28756
rect 19208 28744 19214 28756
rect 19797 28747 19855 28753
rect 19797 28744 19809 28747
rect 19208 28716 19809 28744
rect 19208 28704 19214 28716
rect 19797 28713 19809 28716
rect 19843 28713 19855 28747
rect 19797 28707 19855 28713
rect 19886 28704 19892 28756
rect 19944 28704 19950 28756
rect 19978 28704 19984 28756
rect 20036 28744 20042 28756
rect 21913 28747 21971 28753
rect 20036 28716 20392 28744
rect 20036 28704 20042 28716
rect 19334 28676 19340 28688
rect 18800 28648 19340 28676
rect 18693 28639 18751 28645
rect 17589 28611 17647 28617
rect 17589 28577 17601 28611
rect 17635 28608 17647 28611
rect 18708 28608 18736 28639
rect 19334 28636 19340 28648
rect 19392 28636 19398 28688
rect 19904 28676 19932 28704
rect 19904 28648 20116 28676
rect 19794 28608 19800 28620
rect 17635 28580 18644 28608
rect 18708 28580 19800 28608
rect 17635 28577 17647 28580
rect 17589 28571 17647 28577
rect 15657 28543 15715 28549
rect 15657 28509 15669 28543
rect 15703 28540 15715 28543
rect 16022 28540 16028 28552
rect 15703 28512 16028 28540
rect 15703 28509 15715 28512
rect 15657 28503 15715 28509
rect 16022 28500 16028 28512
rect 16080 28500 16086 28552
rect 16301 28543 16359 28549
rect 16301 28509 16313 28543
rect 16347 28540 16359 28543
rect 16942 28540 16948 28552
rect 16347 28512 16948 28540
rect 16347 28509 16359 28512
rect 16301 28503 16359 28509
rect 16942 28500 16948 28512
rect 17000 28500 17006 28552
rect 17313 28543 17371 28549
rect 17313 28509 17325 28543
rect 17359 28540 17371 28543
rect 18414 28540 18420 28552
rect 17359 28512 18420 28540
rect 17359 28509 17371 28512
rect 17313 28503 17371 28509
rect 18414 28500 18420 28512
rect 18472 28500 18478 28552
rect 16114 28472 16120 28484
rect 16075 28444 16120 28472
rect 16114 28432 16120 28444
rect 16172 28432 16178 28484
rect 16485 28475 16543 28481
rect 16485 28441 16497 28475
rect 16531 28472 16543 28475
rect 17405 28475 17463 28481
rect 17405 28472 17417 28475
rect 16531 28444 17417 28472
rect 16531 28441 16543 28444
rect 16485 28435 16543 28441
rect 17405 28441 17417 28444
rect 17451 28441 17463 28475
rect 18322 28472 18328 28484
rect 18283 28444 18328 28472
rect 17405 28435 17463 28441
rect 18322 28432 18328 28444
rect 18380 28432 18386 28484
rect 18616 28472 18644 28580
rect 19794 28568 19800 28580
rect 19852 28568 19858 28620
rect 20088 28617 20116 28648
rect 20254 28636 20260 28688
rect 20312 28636 20318 28688
rect 20051 28611 20116 28617
rect 20051 28577 20063 28611
rect 20097 28580 20116 28611
rect 20156 28611 20214 28617
rect 20097 28577 20109 28580
rect 20051 28571 20109 28577
rect 20156 28577 20168 28611
rect 20202 28608 20214 28611
rect 20272 28608 20300 28636
rect 20202 28580 20300 28608
rect 20364 28608 20392 28716
rect 21913 28713 21925 28747
rect 21959 28744 21971 28747
rect 22370 28744 22376 28756
rect 21959 28716 22376 28744
rect 21959 28713 21971 28716
rect 21913 28707 21971 28713
rect 22370 28704 22376 28716
rect 22428 28704 22434 28756
rect 23842 28744 23848 28756
rect 23803 28716 23848 28744
rect 23842 28704 23848 28716
rect 23900 28704 23906 28756
rect 24949 28747 25007 28753
rect 24949 28744 24961 28747
rect 24796 28716 24961 28744
rect 20438 28636 20444 28688
rect 20496 28676 20502 28688
rect 20993 28679 21051 28685
rect 20993 28676 21005 28679
rect 20496 28648 21005 28676
rect 20496 28636 20502 28648
rect 20993 28645 21005 28648
rect 21039 28645 21051 28679
rect 20993 28639 21051 28645
rect 23658 28636 23664 28688
rect 23716 28676 23722 28688
rect 24796 28676 24824 28716
rect 24949 28713 24961 28716
rect 24995 28744 25007 28747
rect 27154 28744 27160 28756
rect 24995 28716 27160 28744
rect 24995 28713 25007 28716
rect 24949 28707 25007 28713
rect 27154 28704 27160 28716
rect 27212 28704 27218 28756
rect 27614 28704 27620 28756
rect 27672 28744 27678 28756
rect 27709 28747 27767 28753
rect 27709 28744 27721 28747
rect 27672 28716 27721 28744
rect 27672 28704 27678 28716
rect 27709 28713 27721 28716
rect 27755 28713 27767 28747
rect 30374 28744 30380 28756
rect 27709 28707 27767 28713
rect 28460 28716 30380 28744
rect 27522 28676 27528 28688
rect 23716 28648 24824 28676
rect 24872 28648 27528 28676
rect 23716 28636 23722 28648
rect 20364 28580 21036 28608
rect 20202 28577 20214 28580
rect 20156 28571 20214 28577
rect 19426 28500 19432 28552
rect 19484 28540 19490 28552
rect 19702 28540 19708 28552
rect 19484 28512 19708 28540
rect 19484 28500 19490 28512
rect 19702 28500 19708 28512
rect 19760 28540 19766 28552
rect 19955 28543 20013 28549
rect 19955 28540 19967 28543
rect 19760 28512 19967 28540
rect 19760 28500 19766 28512
rect 19955 28509 19967 28512
rect 20001 28509 20013 28543
rect 19955 28503 20013 28509
rect 20250 28543 20308 28549
rect 20250 28509 20262 28543
rect 20296 28509 20308 28543
rect 20250 28503 20308 28509
rect 19794 28472 19800 28484
rect 18616 28444 19800 28472
rect 19794 28432 19800 28444
rect 19852 28432 19858 28484
rect 20272 28472 20300 28503
rect 20438 28500 20444 28552
rect 20496 28540 20502 28552
rect 20622 28540 20628 28552
rect 20496 28512 20628 28540
rect 20496 28500 20502 28512
rect 20622 28500 20628 28512
rect 20680 28500 20686 28552
rect 20714 28500 20720 28552
rect 20772 28540 20778 28552
rect 21008 28549 21036 28580
rect 20809 28543 20867 28549
rect 20809 28540 20821 28543
rect 20772 28512 20821 28540
rect 20772 28500 20778 28512
rect 20809 28509 20821 28512
rect 20855 28509 20867 28543
rect 20809 28503 20867 28509
rect 20993 28543 21051 28549
rect 20993 28509 21005 28543
rect 21039 28509 21051 28543
rect 21818 28540 21824 28552
rect 20993 28503 21051 28509
rect 21100 28512 21824 28540
rect 21100 28472 21128 28512
rect 21818 28500 21824 28512
rect 21876 28500 21882 28552
rect 22002 28540 22008 28552
rect 21963 28512 22008 28540
rect 22002 28500 22008 28512
rect 22060 28500 22066 28552
rect 22646 28500 22652 28552
rect 22704 28540 22710 28552
rect 24872 28549 24900 28648
rect 27522 28636 27528 28648
rect 27580 28636 27586 28688
rect 27798 28568 27804 28620
rect 27856 28608 27862 28620
rect 28460 28617 28488 28716
rect 30374 28704 30380 28716
rect 30432 28744 30438 28756
rect 31018 28744 31024 28756
rect 30432 28716 31024 28744
rect 30432 28704 30438 28716
rect 31018 28704 31024 28716
rect 31076 28704 31082 28756
rect 31941 28747 31999 28753
rect 31941 28713 31953 28747
rect 31987 28744 31999 28747
rect 33778 28744 33784 28756
rect 31987 28716 33784 28744
rect 31987 28713 31999 28716
rect 31941 28707 31999 28713
rect 33778 28704 33784 28716
rect 33836 28704 33842 28756
rect 34885 28747 34943 28753
rect 34885 28713 34897 28747
rect 34931 28744 34943 28747
rect 35526 28744 35532 28756
rect 34931 28716 35532 28744
rect 34931 28713 34943 28716
rect 34885 28707 34943 28713
rect 35526 28704 35532 28716
rect 35584 28704 35590 28756
rect 36817 28747 36875 28753
rect 36817 28713 36829 28747
rect 36863 28744 36875 28747
rect 37274 28744 37280 28756
rect 36863 28716 37280 28744
rect 36863 28713 36875 28716
rect 36817 28707 36875 28713
rect 37274 28704 37280 28716
rect 37332 28744 37338 28756
rect 37642 28744 37648 28756
rect 37332 28716 37648 28744
rect 37332 28704 37338 28716
rect 37642 28704 37648 28716
rect 37700 28744 37706 28756
rect 37921 28747 37979 28753
rect 37921 28744 37933 28747
rect 37700 28716 37933 28744
rect 37700 28704 37706 28716
rect 37921 28713 37933 28716
rect 37967 28713 37979 28747
rect 37921 28707 37979 28713
rect 30558 28636 30564 28688
rect 30616 28676 30622 28688
rect 32214 28676 32220 28688
rect 30616 28648 32220 28676
rect 30616 28636 30622 28648
rect 32214 28636 32220 28648
rect 32272 28676 32278 28688
rect 34330 28676 34336 28688
rect 32272 28648 33364 28676
rect 32272 28636 32278 28648
rect 28445 28611 28503 28617
rect 28445 28608 28457 28611
rect 27856 28580 28457 28608
rect 27856 28568 27862 28580
rect 28445 28577 28457 28580
rect 28491 28577 28503 28611
rect 28445 28571 28503 28577
rect 28718 28568 28724 28620
rect 28776 28608 28782 28620
rect 31478 28608 31484 28620
rect 28776 28580 31484 28608
rect 28776 28568 28782 28580
rect 31478 28568 31484 28580
rect 31536 28568 31542 28620
rect 31846 28568 31852 28620
rect 31904 28608 31910 28620
rect 31904 28580 32812 28608
rect 31904 28568 31910 28580
rect 22833 28543 22891 28549
rect 22833 28540 22845 28543
rect 22704 28512 22845 28540
rect 22704 28500 22710 28512
rect 22833 28509 22845 28512
rect 22879 28509 22891 28543
rect 22833 28503 22891 28509
rect 23017 28543 23075 28549
rect 23017 28509 23029 28543
rect 23063 28540 23075 28543
rect 24857 28543 24915 28549
rect 24857 28540 24869 28543
rect 23063 28512 24869 28540
rect 23063 28509 23075 28512
rect 23017 28503 23075 28509
rect 24857 28509 24869 28512
rect 24903 28509 24915 28543
rect 24857 28503 24915 28509
rect 25866 28500 25872 28552
rect 25924 28540 25930 28552
rect 26053 28543 26111 28549
rect 26053 28540 26065 28543
rect 25924 28512 26065 28540
rect 25924 28500 25930 28512
rect 26053 28509 26065 28512
rect 26099 28509 26111 28543
rect 26053 28503 26111 28509
rect 26329 28543 26387 28549
rect 26329 28509 26341 28543
rect 26375 28540 26387 28543
rect 26970 28540 26976 28552
rect 26375 28512 26976 28540
rect 26375 28509 26387 28512
rect 26329 28503 26387 28509
rect 20272 28444 21128 28472
rect 21361 28475 21419 28481
rect 21361 28441 21373 28475
rect 21407 28441 21419 28475
rect 23474 28472 23480 28484
rect 23387 28444 23480 28472
rect 21361 28435 21419 28441
rect 18535 28407 18593 28413
rect 18535 28373 18547 28407
rect 18581 28404 18593 28407
rect 18966 28404 18972 28416
rect 18581 28376 18972 28404
rect 18581 28373 18593 28376
rect 18535 28367 18593 28373
rect 18966 28364 18972 28376
rect 19024 28364 19030 28416
rect 19978 28364 19984 28416
rect 20036 28404 20042 28416
rect 21376 28404 21404 28435
rect 23474 28432 23480 28444
rect 23532 28432 23538 28484
rect 23566 28432 23572 28484
rect 23624 28472 23630 28484
rect 23661 28475 23719 28481
rect 23661 28472 23673 28475
rect 23624 28444 23673 28472
rect 23624 28432 23630 28444
rect 23661 28441 23673 28444
rect 23707 28472 23719 28475
rect 23934 28472 23940 28484
rect 23707 28444 23940 28472
rect 23707 28441 23719 28444
rect 23661 28435 23719 28441
rect 23934 28432 23940 28444
rect 23992 28472 23998 28484
rect 26344 28472 26372 28503
rect 26970 28500 26976 28512
rect 27028 28500 27034 28552
rect 27154 28500 27160 28552
rect 27212 28549 27218 28552
rect 27212 28543 27235 28549
rect 27223 28509 27235 28543
rect 27525 28543 27583 28549
rect 27525 28540 27537 28543
rect 27212 28503 27235 28509
rect 27264 28512 27537 28540
rect 27212 28500 27218 28503
rect 23992 28444 26372 28472
rect 26421 28475 26479 28481
rect 23992 28432 23998 28444
rect 26421 28441 26433 28475
rect 26467 28472 26479 28475
rect 27062 28472 27068 28484
rect 26467 28444 27068 28472
rect 26467 28441 26479 28444
rect 26421 28435 26479 28441
rect 20036 28376 21404 28404
rect 20036 28364 20042 28376
rect 22002 28364 22008 28416
rect 22060 28404 22066 28416
rect 23382 28404 23388 28416
rect 22060 28376 23388 28404
rect 22060 28364 22066 28376
rect 23382 28364 23388 28376
rect 23440 28364 23446 28416
rect 23492 28404 23520 28432
rect 23750 28404 23756 28416
rect 23492 28376 23756 28404
rect 23750 28364 23756 28376
rect 23808 28364 23814 28416
rect 24762 28364 24768 28416
rect 24820 28404 24826 28416
rect 26436 28404 26464 28435
rect 27062 28432 27068 28444
rect 27120 28432 27126 28484
rect 27264 28416 27292 28512
rect 27525 28509 27537 28512
rect 27571 28509 27583 28543
rect 28166 28540 28172 28552
rect 28127 28512 28172 28540
rect 27525 28503 27583 28509
rect 28166 28500 28172 28512
rect 28224 28500 28230 28552
rect 29454 28500 29460 28552
rect 29512 28500 29518 28552
rect 30374 28500 30380 28552
rect 30432 28540 30438 28552
rect 30837 28543 30895 28549
rect 30837 28540 30849 28543
rect 30432 28512 30849 28540
rect 30432 28500 30438 28512
rect 30837 28509 30849 28512
rect 30883 28509 30895 28543
rect 31018 28540 31024 28552
rect 30979 28512 31024 28540
rect 30837 28503 30895 28509
rect 31018 28500 31024 28512
rect 31076 28500 31082 28552
rect 32030 28500 32036 28552
rect 32088 28540 32094 28552
rect 32125 28543 32183 28549
rect 32125 28540 32137 28543
rect 32088 28512 32137 28540
rect 32088 28500 32094 28512
rect 32125 28509 32137 28512
rect 32171 28509 32183 28543
rect 32125 28503 32183 28509
rect 32214 28500 32220 28552
rect 32272 28540 32278 28552
rect 32677 28543 32735 28549
rect 32677 28540 32689 28543
rect 32272 28512 32689 28540
rect 32272 28500 32278 28512
rect 32677 28509 32689 28512
rect 32723 28509 32735 28543
rect 32677 28503 32735 28509
rect 32784 28534 32812 28580
rect 33336 28549 33364 28648
rect 33520 28648 34336 28676
rect 33410 28568 33416 28620
rect 33468 28608 33474 28620
rect 33520 28608 33548 28648
rect 34330 28636 34336 28648
rect 34388 28636 34394 28688
rect 34698 28636 34704 28688
rect 34756 28676 34762 28688
rect 35544 28676 35572 28704
rect 34756 28648 35020 28676
rect 35544 28648 37228 28676
rect 34756 28636 34762 28648
rect 33468 28580 33548 28608
rect 33468 28568 33474 28580
rect 33520 28549 33548 28580
rect 34057 28611 34115 28617
rect 34057 28577 34069 28611
rect 34103 28608 34115 28611
rect 34790 28608 34796 28620
rect 34103 28580 34796 28608
rect 34103 28577 34115 28580
rect 34057 28571 34115 28577
rect 34790 28568 34796 28580
rect 34848 28568 34854 28620
rect 34992 28617 35020 28648
rect 34977 28611 35035 28617
rect 34977 28577 34989 28611
rect 35023 28577 35035 28611
rect 34977 28571 35035 28577
rect 32861 28543 32919 28549
rect 32861 28534 32873 28543
rect 32784 28509 32873 28534
rect 32907 28509 32919 28543
rect 32784 28506 32919 28509
rect 32861 28503 32919 28506
rect 33321 28543 33379 28549
rect 33321 28509 33333 28543
rect 33367 28509 33379 28543
rect 33321 28503 33379 28509
rect 33505 28543 33563 28549
rect 33505 28509 33517 28543
rect 33551 28509 33563 28543
rect 33962 28540 33968 28552
rect 33923 28512 33968 28540
rect 33505 28503 33563 28509
rect 33962 28500 33968 28512
rect 34020 28500 34026 28552
rect 34149 28543 34207 28549
rect 34149 28509 34161 28543
rect 34195 28509 34207 28543
rect 34149 28503 34207 28509
rect 27341 28475 27399 28481
rect 27341 28441 27353 28475
rect 27387 28441 27399 28475
rect 27341 28435 27399 28441
rect 27433 28475 27491 28481
rect 27433 28441 27445 28475
rect 27479 28472 27491 28475
rect 28534 28472 28540 28484
rect 27479 28444 28540 28472
rect 27479 28441 27491 28444
rect 27433 28435 27491 28441
rect 24820 28376 26464 28404
rect 24820 28364 24826 28376
rect 27246 28364 27252 28416
rect 27304 28364 27310 28416
rect 27356 28404 27384 28435
rect 28534 28432 28540 28444
rect 28592 28432 28598 28484
rect 29472 28472 29500 28500
rect 30009 28475 30067 28481
rect 30009 28472 30021 28475
rect 29472 28444 30021 28472
rect 30009 28441 30021 28444
rect 30055 28472 30067 28475
rect 31846 28472 31852 28484
rect 30055 28444 31852 28472
rect 30055 28441 30067 28444
rect 30009 28435 30067 28441
rect 31846 28432 31852 28444
rect 31904 28432 31910 28484
rect 31941 28475 31999 28481
rect 31941 28441 31953 28475
rect 31987 28472 31999 28475
rect 32306 28472 32312 28484
rect 31987 28444 32312 28472
rect 31987 28441 31999 28444
rect 31941 28435 31999 28441
rect 32306 28432 32312 28444
rect 32364 28432 32370 28484
rect 33413 28475 33471 28481
rect 32416 28444 32904 28472
rect 27982 28404 27988 28416
rect 27356 28376 27988 28404
rect 27982 28364 27988 28376
rect 28040 28404 28046 28416
rect 30101 28407 30159 28413
rect 30101 28404 30113 28407
rect 28040 28376 30113 28404
rect 28040 28364 28046 28376
rect 30101 28373 30113 28376
rect 30147 28373 30159 28407
rect 30101 28367 30159 28373
rect 30190 28364 30196 28416
rect 30248 28404 30254 28416
rect 30929 28407 30987 28413
rect 30929 28404 30941 28407
rect 30248 28376 30941 28404
rect 30248 28364 30254 28376
rect 30929 28373 30941 28376
rect 30975 28373 30987 28407
rect 30929 28367 30987 28373
rect 32214 28364 32220 28416
rect 32272 28404 32278 28416
rect 32416 28404 32444 28444
rect 32272 28376 32444 28404
rect 32272 28364 32278 28376
rect 32674 28364 32680 28416
rect 32732 28404 32738 28416
rect 32769 28407 32827 28413
rect 32769 28404 32781 28407
rect 32732 28376 32781 28404
rect 32732 28364 32738 28376
rect 32769 28373 32781 28376
rect 32815 28373 32827 28407
rect 32876 28404 32904 28444
rect 33413 28441 33425 28475
rect 33459 28472 33471 28475
rect 33870 28472 33876 28484
rect 33459 28444 33876 28472
rect 33459 28441 33471 28444
rect 33413 28435 33471 28441
rect 33870 28432 33876 28444
rect 33928 28472 33934 28484
rect 34164 28472 34192 28503
rect 34514 28500 34520 28552
rect 34572 28540 34578 28552
rect 34701 28543 34759 28549
rect 34701 28540 34713 28543
rect 34572 28512 34713 28540
rect 34572 28500 34578 28512
rect 34701 28509 34713 28512
rect 34747 28509 34759 28543
rect 34701 28503 34759 28509
rect 35805 28543 35863 28549
rect 35805 28509 35817 28543
rect 35851 28540 35863 28543
rect 35894 28540 35900 28552
rect 35851 28512 35900 28540
rect 35851 28509 35863 28512
rect 35805 28503 35863 28509
rect 35894 28500 35900 28512
rect 35952 28500 35958 28552
rect 36538 28500 36544 28552
rect 36596 28540 36602 28552
rect 37200 28549 37228 28648
rect 37001 28543 37059 28549
rect 37001 28540 37013 28543
rect 36596 28512 37013 28540
rect 36596 28500 36602 28512
rect 37001 28509 37013 28512
rect 37047 28509 37059 28543
rect 37001 28503 37059 28509
rect 37185 28543 37243 28549
rect 37185 28509 37197 28543
rect 37231 28509 37243 28543
rect 37185 28503 37243 28509
rect 37274 28500 37280 28552
rect 37332 28540 37338 28552
rect 37332 28512 37377 28540
rect 37332 28500 37338 28512
rect 35986 28472 35992 28484
rect 33928 28444 34192 28472
rect 35947 28444 35992 28472
rect 33928 28432 33934 28444
rect 35986 28432 35992 28444
rect 36044 28432 36050 28484
rect 36096 28444 36676 28472
rect 36096 28404 36124 28444
rect 32876 28376 36124 28404
rect 36173 28407 36231 28413
rect 32769 28367 32827 28373
rect 36173 28373 36185 28407
rect 36219 28404 36231 28407
rect 36538 28404 36544 28416
rect 36219 28376 36544 28404
rect 36219 28373 36231 28376
rect 36173 28367 36231 28373
rect 36538 28364 36544 28376
rect 36596 28364 36602 28416
rect 36648 28404 36676 28444
rect 37458 28432 37464 28484
rect 37516 28472 37522 28484
rect 37737 28475 37795 28481
rect 37737 28472 37749 28475
rect 37516 28444 37749 28472
rect 37516 28432 37522 28444
rect 37737 28441 37749 28444
rect 37783 28441 37795 28475
rect 37737 28435 37795 28441
rect 37918 28432 37924 28484
rect 37976 28481 37982 28484
rect 37976 28475 37995 28481
rect 37983 28441 37995 28475
rect 37976 28435 37995 28441
rect 37976 28432 37982 28435
rect 37366 28404 37372 28416
rect 36648 28376 37372 28404
rect 37366 28364 37372 28376
rect 37424 28364 37430 28416
rect 38102 28404 38108 28416
rect 38063 28376 38108 28404
rect 38102 28364 38108 28376
rect 38160 28364 38166 28416
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 16114 28160 16120 28212
rect 16172 28200 16178 28212
rect 17313 28203 17371 28209
rect 17313 28200 17325 28203
rect 16172 28172 17325 28200
rect 16172 28160 16178 28172
rect 17313 28169 17325 28172
rect 17359 28169 17371 28203
rect 17313 28163 17371 28169
rect 18230 28160 18236 28212
rect 18288 28200 18294 28212
rect 18509 28203 18567 28209
rect 18509 28200 18521 28203
rect 18288 28172 18521 28200
rect 18288 28160 18294 28172
rect 18509 28169 18521 28172
rect 18555 28169 18567 28203
rect 18509 28163 18567 28169
rect 18800 28172 19840 28200
rect 16945 28135 17003 28141
rect 16945 28101 16957 28135
rect 16991 28132 17003 28135
rect 17034 28132 17040 28144
rect 16991 28104 17040 28132
rect 16991 28101 17003 28104
rect 16945 28095 17003 28101
rect 17034 28092 17040 28104
rect 17092 28092 17098 28144
rect 17126 28092 17132 28144
rect 17184 28141 17190 28144
rect 17184 28135 17219 28141
rect 17207 28132 17219 28135
rect 17207 28104 17816 28132
rect 17207 28101 17219 28104
rect 17184 28095 17219 28101
rect 17184 28092 17190 28095
rect 13814 28024 13820 28076
rect 13872 28064 13878 28076
rect 15105 28067 15163 28073
rect 15105 28064 15117 28067
rect 13872 28036 15117 28064
rect 13872 28024 13878 28036
rect 15105 28033 15117 28036
rect 15151 28033 15163 28067
rect 15105 28027 15163 28033
rect 14274 27956 14280 28008
rect 14332 27996 14338 28008
rect 14829 27999 14887 28005
rect 14829 27996 14841 27999
rect 14332 27968 14841 27996
rect 14332 27956 14338 27968
rect 14829 27965 14841 27968
rect 14875 27965 14887 27999
rect 17788 27996 17816 28104
rect 17865 28067 17923 28073
rect 17865 28033 17877 28067
rect 17911 28064 17923 28067
rect 18322 28064 18328 28076
rect 17911 28036 18328 28064
rect 17911 28033 17923 28036
rect 17865 28027 17923 28033
rect 18322 28024 18328 28036
rect 18380 28064 18386 28076
rect 18693 28067 18751 28073
rect 18693 28064 18705 28067
rect 18380 28036 18705 28064
rect 18380 28024 18386 28036
rect 18693 28033 18705 28036
rect 18739 28064 18751 28067
rect 18800 28064 18828 28172
rect 18877 28135 18935 28141
rect 18877 28101 18889 28135
rect 18923 28132 18935 28135
rect 19334 28132 19340 28144
rect 18923 28104 19340 28132
rect 18923 28101 18935 28104
rect 18877 28095 18935 28101
rect 19334 28092 19340 28104
rect 19392 28132 19398 28144
rect 19812 28132 19840 28172
rect 20622 28160 20628 28212
rect 20680 28160 20686 28212
rect 23385 28203 23443 28209
rect 23385 28169 23397 28203
rect 23431 28200 23443 28203
rect 24946 28200 24952 28212
rect 23431 28172 24952 28200
rect 23431 28169 23443 28172
rect 23385 28163 23443 28169
rect 24946 28160 24952 28172
rect 25004 28160 25010 28212
rect 25038 28160 25044 28212
rect 25096 28200 25102 28212
rect 25958 28200 25964 28212
rect 25096 28172 25964 28200
rect 25096 28160 25102 28172
rect 25958 28160 25964 28172
rect 26016 28200 26022 28212
rect 26016 28172 27568 28200
rect 26016 28160 26022 28172
rect 20640 28132 20668 28160
rect 19392 28104 19748 28132
rect 19392 28092 19398 28104
rect 18739 28036 18828 28064
rect 18739 28033 18751 28036
rect 18693 28027 18751 28033
rect 18966 28024 18972 28076
rect 19024 28064 19030 28076
rect 19024 28036 19656 28064
rect 19024 28024 19030 28036
rect 19426 27996 19432 28008
rect 17788 27968 18828 27996
rect 19387 27968 19432 27996
rect 14829 27959 14887 27965
rect 15841 27863 15899 27869
rect 15841 27829 15853 27863
rect 15887 27860 15899 27863
rect 16850 27860 16856 27872
rect 15887 27832 16856 27860
rect 15887 27829 15899 27832
rect 15841 27823 15899 27829
rect 16850 27820 16856 27832
rect 16908 27820 16914 27872
rect 17129 27863 17187 27869
rect 17129 27829 17141 27863
rect 17175 27860 17187 27863
rect 17218 27860 17224 27872
rect 17175 27832 17224 27860
rect 17175 27829 17187 27832
rect 17129 27823 17187 27829
rect 17218 27820 17224 27832
rect 17276 27820 17282 27872
rect 17957 27863 18015 27869
rect 17957 27829 17969 27863
rect 18003 27860 18015 27863
rect 18690 27860 18696 27872
rect 18003 27832 18696 27860
rect 18003 27829 18015 27832
rect 17957 27823 18015 27829
rect 18690 27820 18696 27832
rect 18748 27820 18754 27872
rect 18800 27860 18828 27968
rect 19426 27956 19432 27968
rect 19484 27956 19490 28008
rect 19628 28005 19656 28036
rect 19720 28008 19748 28104
rect 19812 28104 20668 28132
rect 20809 28135 20867 28141
rect 19812 28073 19840 28104
rect 20809 28101 20821 28135
rect 20855 28132 20867 28135
rect 20855 28104 20944 28132
rect 20855 28101 20867 28104
rect 20809 28095 20867 28101
rect 19797 28067 19855 28073
rect 19797 28033 19809 28067
rect 19843 28033 19855 28067
rect 19797 28027 19855 28033
rect 19889 28067 19947 28073
rect 19889 28033 19901 28067
rect 19935 28064 19947 28067
rect 19978 28064 19984 28076
rect 19935 28036 19984 28064
rect 19935 28033 19947 28036
rect 19889 28027 19947 28033
rect 19978 28024 19984 28036
rect 20036 28024 20042 28076
rect 20622 28064 20628 28076
rect 20583 28036 20628 28064
rect 20622 28024 20628 28036
rect 20680 28024 20686 28076
rect 20714 28024 20720 28076
rect 20772 28064 20778 28076
rect 20772 28036 20817 28064
rect 20772 28024 20778 28036
rect 19613 27999 19671 28005
rect 19613 27965 19625 27999
rect 19659 27965 19671 27999
rect 19613 27959 19671 27965
rect 19628 27928 19656 27959
rect 19702 27956 19708 28008
rect 19760 27996 19766 28008
rect 19760 27968 19805 27996
rect 19760 27956 19766 27968
rect 20254 27956 20260 28008
rect 20312 27996 20318 28008
rect 20916 27996 20944 28104
rect 23014 28092 23020 28144
rect 23072 28132 23078 28144
rect 27540 28132 27568 28172
rect 28166 28160 28172 28212
rect 28224 28200 28230 28212
rect 28445 28203 28503 28209
rect 28445 28200 28457 28203
rect 28224 28172 28457 28200
rect 28224 28160 28230 28172
rect 28445 28169 28457 28172
rect 28491 28200 28503 28203
rect 29546 28200 29552 28212
rect 28491 28172 29552 28200
rect 28491 28169 28503 28172
rect 28445 28163 28503 28169
rect 29546 28160 29552 28172
rect 29604 28160 29610 28212
rect 30101 28203 30159 28209
rect 30101 28169 30113 28203
rect 30147 28200 30159 28203
rect 30926 28200 30932 28212
rect 30147 28172 30932 28200
rect 30147 28169 30159 28172
rect 30101 28163 30159 28169
rect 30926 28160 30932 28172
rect 30984 28160 30990 28212
rect 31389 28203 31447 28209
rect 31389 28169 31401 28203
rect 31435 28169 31447 28203
rect 31389 28163 31447 28169
rect 28718 28132 28724 28144
rect 23072 28104 27476 28132
rect 27540 28104 28724 28132
rect 23072 28092 23078 28104
rect 20993 28067 21051 28073
rect 20993 28042 21005 28067
rect 21039 28042 21051 28067
rect 21085 28067 21143 28073
rect 20312 27968 20944 27996
rect 20990 27990 20996 28042
rect 21048 27990 21054 28042
rect 21085 28033 21097 28067
rect 21131 28033 21143 28067
rect 21085 28027 21143 28033
rect 21100 27996 21128 28027
rect 21174 28024 21180 28076
rect 21232 28064 21238 28076
rect 21821 28067 21879 28073
rect 21821 28064 21833 28067
rect 21232 28036 21833 28064
rect 21232 28024 21238 28036
rect 21821 28033 21833 28036
rect 21867 28033 21879 28067
rect 21821 28027 21879 28033
rect 22094 28024 22100 28076
rect 22152 28064 22158 28076
rect 22557 28067 22615 28073
rect 22557 28064 22569 28067
rect 22152 28036 22569 28064
rect 22152 28024 22158 28036
rect 22557 28033 22569 28036
rect 22603 28033 22615 28067
rect 22557 28027 22615 28033
rect 22738 28024 22744 28076
rect 22796 28064 22802 28076
rect 23201 28067 23259 28073
rect 23201 28064 23213 28067
rect 22796 28036 23213 28064
rect 22796 28024 22802 28036
rect 23201 28033 23213 28036
rect 23247 28033 23259 28067
rect 23201 28027 23259 28033
rect 24029 28067 24087 28073
rect 24029 28033 24041 28067
rect 24075 28064 24087 28067
rect 24210 28064 24216 28076
rect 24075 28036 24216 28064
rect 24075 28033 24087 28036
rect 24029 28027 24087 28033
rect 24210 28024 24216 28036
rect 24268 28024 24274 28076
rect 24762 28064 24768 28076
rect 24723 28036 24768 28064
rect 24762 28024 24768 28036
rect 24820 28024 24826 28076
rect 24949 28067 25007 28073
rect 24949 28033 24961 28067
rect 24995 28064 25007 28067
rect 25038 28064 25044 28076
rect 24995 28036 25044 28064
rect 24995 28033 25007 28036
rect 24949 28027 25007 28033
rect 25038 28024 25044 28036
rect 25096 28024 25102 28076
rect 25222 28024 25228 28076
rect 25280 28064 25286 28076
rect 27448 28073 27476 28104
rect 28718 28092 28724 28104
rect 28776 28092 28782 28144
rect 28810 28092 28816 28144
rect 28868 28132 28874 28144
rect 31110 28132 31116 28144
rect 28868 28104 30972 28132
rect 31071 28104 31116 28132
rect 28868 28092 28874 28104
rect 25777 28067 25835 28073
rect 25777 28064 25789 28067
rect 25280 28036 25789 28064
rect 25280 28024 25286 28036
rect 25777 28033 25789 28036
rect 25823 28033 25835 28067
rect 25777 28027 25835 28033
rect 25961 28067 26019 28073
rect 25961 28033 25973 28067
rect 26007 28033 26019 28067
rect 25961 28027 26019 28033
rect 27433 28067 27491 28073
rect 27433 28033 27445 28067
rect 27479 28033 27491 28067
rect 27433 28027 27491 28033
rect 21266 27996 21272 28008
rect 21100 27968 21272 27996
rect 20312 27956 20318 27968
rect 21266 27956 21272 27968
rect 21324 27956 21330 28008
rect 23750 27956 23756 28008
rect 23808 27996 23814 28008
rect 25976 27996 26004 28027
rect 23808 27968 26004 27996
rect 27448 27996 27476 28027
rect 27706 28024 27712 28076
rect 27764 28064 27770 28076
rect 28166 28064 28172 28076
rect 27764 28036 28172 28064
rect 27764 28024 27770 28036
rect 28166 28024 28172 28036
rect 28224 28024 28230 28076
rect 28353 28067 28411 28073
rect 28353 28033 28365 28067
rect 28399 28064 28411 28067
rect 28902 28064 28908 28076
rect 28399 28036 28908 28064
rect 28399 28033 28411 28036
rect 28353 28027 28411 28033
rect 28902 28024 28908 28036
rect 28960 28024 28966 28076
rect 29104 28073 29132 28104
rect 30944 28076 30972 28104
rect 31110 28092 31116 28104
rect 31168 28092 31174 28144
rect 31404 28132 31432 28163
rect 31478 28160 31484 28212
rect 31536 28200 31542 28212
rect 31536 28172 34376 28200
rect 31536 28160 31542 28172
rect 31846 28132 31852 28144
rect 31404 28104 31852 28132
rect 31846 28092 31852 28104
rect 31904 28132 31910 28144
rect 32398 28132 32404 28144
rect 31904 28104 32260 28132
rect 32311 28104 32404 28132
rect 31904 28092 31910 28104
rect 29089 28067 29147 28073
rect 29089 28033 29101 28067
rect 29135 28033 29147 28067
rect 29089 28027 29147 28033
rect 29178 28024 29184 28076
rect 29236 28064 29242 28076
rect 29273 28067 29331 28073
rect 29273 28064 29285 28067
rect 29236 28036 29285 28064
rect 29236 28024 29242 28036
rect 29273 28033 29285 28036
rect 29319 28033 29331 28067
rect 29273 28027 29331 28033
rect 28074 27996 28080 28008
rect 27448 27968 28080 27996
rect 23808 27956 23814 27968
rect 28074 27956 28080 27968
rect 28132 27956 28138 28008
rect 29288 27996 29316 28027
rect 29362 28024 29368 28076
rect 29420 28064 29426 28076
rect 29730 28064 29736 28076
rect 29420 28036 29736 28064
rect 29420 28024 29426 28036
rect 29730 28024 29736 28036
rect 29788 28064 29794 28076
rect 29825 28067 29883 28073
rect 29825 28064 29837 28067
rect 29788 28036 29837 28064
rect 29788 28024 29794 28036
rect 29825 28033 29837 28036
rect 29871 28033 29883 28067
rect 30834 28064 30840 28076
rect 29825 28027 29883 28033
rect 30024 28036 30840 28064
rect 29638 27996 29644 28008
rect 29288 27968 29644 27996
rect 29638 27956 29644 27968
rect 29696 27956 29702 28008
rect 30024 27996 30052 28036
rect 30834 28024 30840 28036
rect 30892 28024 30898 28076
rect 30926 28024 30932 28076
rect 30984 28064 30990 28076
rect 31021 28067 31079 28073
rect 31021 28064 31033 28067
rect 30984 28036 31033 28064
rect 30984 28024 30990 28036
rect 31021 28033 31033 28036
rect 31067 28033 31079 28067
rect 31021 28027 31079 28033
rect 31205 28067 31263 28073
rect 31205 28033 31217 28067
rect 31251 28064 31263 28067
rect 31251 28036 31432 28064
rect 31251 28033 31263 28036
rect 31205 28027 31263 28033
rect 31404 28008 31432 28036
rect 31938 28024 31944 28076
rect 31996 28064 32002 28076
rect 32232 28073 32260 28104
rect 32398 28092 32404 28104
rect 32456 28132 32462 28144
rect 32456 28104 33088 28132
rect 32456 28092 32462 28104
rect 32125 28067 32183 28073
rect 32125 28064 32137 28067
rect 31996 28036 32137 28064
rect 31996 28024 32002 28036
rect 32125 28033 32137 28036
rect 32171 28033 32183 28067
rect 32125 28027 32183 28033
rect 32217 28067 32275 28073
rect 32217 28033 32229 28067
rect 32263 28033 32275 28067
rect 32217 28027 32275 28033
rect 32493 28067 32551 28073
rect 32493 28033 32505 28067
rect 32539 28033 32551 28067
rect 32493 28027 32551 28033
rect 32585 28067 32643 28073
rect 32585 28033 32597 28067
rect 32631 28064 32643 28067
rect 32766 28064 32772 28076
rect 32631 28036 32772 28064
rect 32631 28033 32643 28036
rect 32585 28027 32643 28033
rect 29866 27968 30052 27996
rect 20441 27931 20499 27937
rect 20441 27928 20453 27931
rect 19628 27900 20453 27928
rect 20441 27897 20453 27900
rect 20487 27897 20499 27931
rect 22370 27928 22376 27940
rect 20441 27891 20499 27897
rect 20548 27900 22376 27928
rect 20548 27860 20576 27900
rect 22370 27888 22376 27900
rect 22428 27888 22434 27940
rect 22741 27931 22799 27937
rect 22741 27897 22753 27931
rect 22787 27928 22799 27931
rect 26602 27928 26608 27940
rect 22787 27900 26608 27928
rect 22787 27897 22799 27900
rect 22741 27891 22799 27897
rect 26602 27888 26608 27900
rect 26660 27888 26666 27940
rect 27614 27928 27620 27940
rect 27575 27900 27620 27928
rect 27614 27888 27620 27900
rect 27672 27928 27678 27940
rect 29866 27928 29894 27968
rect 30098 27956 30104 28008
rect 30156 27996 30162 28008
rect 30156 27968 30201 27996
rect 30156 27956 30162 27968
rect 30282 27956 30288 28008
rect 30340 27996 30346 28008
rect 31386 27996 31392 28008
rect 30340 27968 31392 27996
rect 30340 27956 30346 27968
rect 31386 27956 31392 27968
rect 31444 27956 31450 28008
rect 32030 27928 32036 27940
rect 27672 27900 29894 27928
rect 30300 27900 32036 27928
rect 27672 27888 27678 27900
rect 18800 27832 20576 27860
rect 21818 27820 21824 27872
rect 21876 27860 21882 27872
rect 21913 27863 21971 27869
rect 21913 27860 21925 27863
rect 21876 27832 21925 27860
rect 21876 27820 21882 27832
rect 21913 27829 21925 27832
rect 21959 27860 21971 27863
rect 22278 27860 22284 27872
rect 21959 27832 22284 27860
rect 21959 27829 21971 27832
rect 21913 27823 21971 27829
rect 22278 27820 22284 27832
rect 22336 27820 22342 27872
rect 24121 27863 24179 27869
rect 24121 27829 24133 27863
rect 24167 27860 24179 27863
rect 25774 27860 25780 27872
rect 24167 27832 25780 27860
rect 24167 27829 24179 27832
rect 24121 27823 24179 27829
rect 25774 27820 25780 27832
rect 25832 27820 25838 27872
rect 25869 27863 25927 27869
rect 25869 27829 25881 27863
rect 25915 27860 25927 27863
rect 25958 27860 25964 27872
rect 25915 27832 25964 27860
rect 25915 27829 25927 27832
rect 25869 27823 25927 27829
rect 25958 27820 25964 27832
rect 26016 27860 26022 27872
rect 27430 27860 27436 27872
rect 26016 27832 27436 27860
rect 26016 27820 26022 27832
rect 27430 27820 27436 27832
rect 27488 27820 27494 27872
rect 28442 27820 28448 27872
rect 28500 27860 28506 27872
rect 28994 27860 29000 27872
rect 28500 27832 29000 27860
rect 28500 27820 28506 27832
rect 28994 27820 29000 27832
rect 29052 27820 29058 27872
rect 29638 27820 29644 27872
rect 29696 27860 29702 27872
rect 29917 27863 29975 27869
rect 29917 27860 29929 27863
rect 29696 27832 29929 27860
rect 29696 27820 29702 27832
rect 29917 27829 29929 27832
rect 29963 27860 29975 27863
rect 30300 27860 30328 27900
rect 32030 27888 32036 27900
rect 32088 27888 32094 27940
rect 32125 27931 32183 27937
rect 32125 27897 32137 27931
rect 32171 27928 32183 27931
rect 32398 27928 32404 27940
rect 32171 27900 32404 27928
rect 32171 27897 32183 27900
rect 32125 27891 32183 27897
rect 32398 27888 32404 27900
rect 32456 27888 32462 27940
rect 32508 27928 32536 28027
rect 32766 28024 32772 28036
rect 32824 28024 32830 28076
rect 32674 27928 32680 27940
rect 32508 27900 32680 27928
rect 32674 27888 32680 27900
rect 32732 27888 32738 27940
rect 33060 27928 33088 28104
rect 33594 28092 33600 28144
rect 33652 28132 33658 28144
rect 33873 28135 33931 28141
rect 33873 28132 33885 28135
rect 33652 28104 33885 28132
rect 33652 28092 33658 28104
rect 33873 28101 33885 28104
rect 33919 28101 33931 28135
rect 33873 28095 33931 28101
rect 33686 28064 33692 28076
rect 33647 28036 33692 28064
rect 33686 28024 33692 28036
rect 33744 28024 33750 28076
rect 34348 28073 34376 28172
rect 34422 28160 34428 28212
rect 34480 28200 34486 28212
rect 37642 28200 37648 28212
rect 34480 28172 34525 28200
rect 37603 28172 37648 28200
rect 34480 28160 34486 28172
rect 37642 28160 37648 28172
rect 37700 28160 37706 28212
rect 34333 28067 34391 28073
rect 34333 28033 34345 28067
rect 34379 28033 34391 28067
rect 34514 28064 34520 28076
rect 34475 28036 34520 28064
rect 34333 28027 34391 28033
rect 34514 28024 34520 28036
rect 34572 28024 34578 28076
rect 34977 28067 35035 28073
rect 34977 28033 34989 28067
rect 35023 28033 35035 28067
rect 34977 28027 35035 28033
rect 35161 28067 35219 28073
rect 35161 28033 35173 28067
rect 35207 28064 35219 28067
rect 35434 28064 35440 28076
rect 35207 28036 35440 28064
rect 35207 28033 35219 28036
rect 35161 28027 35219 28033
rect 33962 27956 33968 28008
rect 34020 27996 34026 28008
rect 34992 27996 35020 28027
rect 35434 28024 35440 28036
rect 35492 28024 35498 28076
rect 35894 28064 35900 28076
rect 35855 28036 35900 28064
rect 35894 28024 35900 28036
rect 35952 28024 35958 28076
rect 35986 28024 35992 28076
rect 36044 28064 36050 28076
rect 36081 28067 36139 28073
rect 36081 28064 36093 28067
rect 36044 28036 36093 28064
rect 36044 28024 36050 28036
rect 36081 28033 36093 28036
rect 36127 28033 36139 28067
rect 36538 28064 36544 28076
rect 36499 28036 36544 28064
rect 36081 28027 36139 28033
rect 36538 28024 36544 28036
rect 36596 28024 36602 28076
rect 36725 28067 36783 28073
rect 36725 28033 36737 28067
rect 36771 28064 36783 28067
rect 37274 28064 37280 28076
rect 36771 28036 37280 28064
rect 36771 28033 36783 28036
rect 36725 28027 36783 28033
rect 36630 27996 36636 28008
rect 34020 27968 35020 27996
rect 36004 27968 36636 27996
rect 34020 27956 34026 27968
rect 36004 27937 36032 27968
rect 36630 27956 36636 27968
rect 36688 27996 36694 28008
rect 36740 27996 36768 28027
rect 37274 28024 37280 28036
rect 37332 28024 37338 28076
rect 37458 28064 37464 28076
rect 37419 28036 37464 28064
rect 37458 28024 37464 28036
rect 37516 28024 37522 28076
rect 37737 28067 37795 28073
rect 37737 28033 37749 28067
rect 37783 28064 37795 28067
rect 37918 28064 37924 28076
rect 37783 28036 37924 28064
rect 37783 28033 37795 28036
rect 37737 28027 37795 28033
rect 37918 28024 37924 28036
rect 37976 28024 37982 28076
rect 36688 27968 36768 27996
rect 36688 27956 36694 27968
rect 35989 27931 36047 27937
rect 33060 27900 35020 27928
rect 29963 27832 30328 27860
rect 29963 27829 29975 27832
rect 29917 27823 29975 27829
rect 31938 27820 31944 27872
rect 31996 27860 32002 27872
rect 33042 27860 33048 27872
rect 31996 27832 33048 27860
rect 31996 27820 32002 27832
rect 33042 27820 33048 27832
rect 33100 27860 33106 27872
rect 33870 27860 33876 27872
rect 33100 27832 33876 27860
rect 33100 27820 33106 27832
rect 33870 27820 33876 27832
rect 33928 27820 33934 27872
rect 34992 27869 35020 27900
rect 35989 27897 36001 27931
rect 36035 27897 36047 27931
rect 35989 27891 36047 27897
rect 34977 27863 35035 27869
rect 34977 27829 34989 27863
rect 35023 27829 35035 27863
rect 36630 27860 36636 27872
rect 36591 27832 36636 27860
rect 34977 27823 35035 27829
rect 36630 27820 36636 27832
rect 36688 27820 36694 27872
rect 37461 27863 37519 27869
rect 37461 27829 37473 27863
rect 37507 27860 37519 27863
rect 37734 27860 37740 27872
rect 37507 27832 37740 27860
rect 37507 27829 37519 27832
rect 37461 27823 37519 27829
rect 37734 27820 37740 27832
rect 37792 27820 37798 27872
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 16942 27656 16948 27668
rect 16903 27628 16948 27656
rect 16942 27616 16948 27628
rect 17000 27616 17006 27668
rect 18141 27659 18199 27665
rect 18141 27625 18153 27659
rect 18187 27656 18199 27659
rect 19429 27659 19487 27665
rect 19429 27656 19441 27659
rect 18187 27628 19441 27656
rect 18187 27625 18199 27628
rect 18141 27619 18199 27625
rect 19429 27625 19441 27628
rect 19475 27625 19487 27659
rect 19429 27619 19487 27625
rect 16393 27591 16451 27597
rect 16393 27557 16405 27591
rect 16439 27588 16451 27591
rect 17770 27588 17776 27600
rect 16439 27560 17776 27588
rect 16439 27557 16451 27560
rect 16393 27551 16451 27557
rect 17770 27548 17776 27560
rect 17828 27548 17834 27600
rect 19444 27588 19472 27619
rect 19702 27616 19708 27668
rect 19760 27656 19766 27668
rect 19981 27659 20039 27665
rect 19981 27656 19993 27659
rect 19760 27628 19993 27656
rect 19760 27616 19766 27628
rect 19981 27625 19993 27628
rect 20027 27625 20039 27659
rect 20346 27656 20352 27668
rect 19981 27619 20039 27625
rect 20088 27628 20352 27656
rect 20088 27588 20116 27628
rect 20346 27616 20352 27628
rect 20404 27616 20410 27668
rect 20990 27616 20996 27668
rect 21048 27656 21054 27668
rect 21177 27659 21235 27665
rect 21177 27656 21189 27659
rect 21048 27628 21189 27656
rect 21048 27616 21054 27628
rect 21177 27625 21189 27628
rect 21223 27656 21235 27659
rect 23014 27656 23020 27668
rect 21223 27628 23020 27656
rect 21223 27625 21235 27628
rect 21177 27619 21235 27625
rect 23014 27616 23020 27628
rect 23072 27616 23078 27668
rect 25866 27656 25872 27668
rect 25827 27628 25872 27656
rect 25866 27616 25872 27628
rect 25924 27616 25930 27668
rect 27617 27659 27675 27665
rect 27617 27625 27629 27659
rect 27663 27656 27675 27659
rect 27890 27656 27896 27668
rect 27663 27628 27896 27656
rect 27663 27625 27675 27628
rect 27617 27619 27675 27625
rect 27890 27616 27896 27628
rect 27948 27616 27954 27668
rect 28313 27659 28371 27665
rect 28313 27656 28325 27659
rect 28308 27625 28325 27656
rect 28359 27625 28371 27659
rect 28308 27619 28371 27625
rect 19444 27560 20116 27588
rect 20162 27548 20168 27600
rect 20220 27588 20226 27600
rect 20220 27560 23060 27588
rect 20220 27548 20226 27560
rect 17126 27520 17132 27532
rect 16960 27492 17132 27520
rect 14274 27412 14280 27464
rect 14332 27452 14338 27464
rect 14461 27455 14519 27461
rect 14461 27452 14473 27455
rect 14332 27424 14473 27452
rect 14332 27412 14338 27424
rect 14461 27421 14473 27424
rect 14507 27421 14519 27455
rect 14734 27452 14740 27464
rect 14695 27424 14740 27452
rect 14461 27415 14519 27421
rect 14734 27412 14740 27424
rect 14792 27412 14798 27464
rect 15930 27412 15936 27464
rect 15988 27452 15994 27464
rect 16960 27461 16988 27492
rect 17126 27480 17132 27492
rect 17184 27480 17190 27532
rect 18598 27520 18604 27532
rect 17788 27492 18604 27520
rect 16209 27455 16267 27461
rect 16209 27452 16221 27455
rect 15988 27424 16221 27452
rect 15988 27412 15994 27424
rect 16209 27421 16221 27424
rect 16255 27421 16267 27455
rect 16209 27415 16267 27421
rect 16945 27455 17003 27461
rect 16945 27421 16957 27455
rect 16991 27421 17003 27455
rect 17218 27452 17224 27464
rect 17179 27424 17224 27452
rect 16945 27415 17003 27421
rect 17218 27412 17224 27424
rect 17276 27412 17282 27464
rect 17788 27461 17816 27492
rect 18598 27480 18604 27492
rect 18656 27520 18662 27532
rect 19334 27520 19340 27532
rect 18656 27492 19340 27520
rect 18656 27480 18662 27492
rect 19334 27480 19340 27492
rect 19392 27520 19398 27532
rect 20622 27520 20628 27532
rect 19392 27492 20628 27520
rect 19392 27480 19398 27492
rect 17773 27455 17831 27461
rect 17773 27421 17785 27455
rect 17819 27421 17831 27455
rect 18046 27452 18052 27464
rect 18007 27424 18052 27452
rect 17773 27415 17831 27421
rect 18046 27412 18052 27424
rect 18104 27412 18110 27464
rect 20162 27452 20168 27464
rect 18156 27424 19472 27452
rect 20123 27424 20168 27452
rect 16758 27384 16764 27396
rect 16132 27356 16764 27384
rect 16132 27328 16160 27356
rect 16758 27344 16764 27356
rect 16816 27344 16822 27396
rect 16850 27344 16856 27396
rect 16908 27384 16914 27396
rect 18156 27384 18184 27424
rect 16908 27356 18184 27384
rect 16908 27344 16914 27356
rect 19242 27344 19248 27396
rect 19300 27384 19306 27396
rect 19337 27387 19395 27393
rect 19337 27384 19349 27387
rect 19300 27356 19349 27384
rect 19300 27344 19306 27356
rect 19337 27353 19349 27356
rect 19383 27353 19395 27387
rect 19444 27384 19472 27424
rect 20162 27412 20168 27424
rect 20220 27412 20226 27464
rect 20456 27461 20484 27492
rect 20622 27480 20628 27492
rect 20680 27480 20686 27532
rect 23032 27529 23060 27560
rect 24762 27548 24768 27600
rect 24820 27588 24826 27600
rect 28074 27588 28080 27600
rect 24820 27560 28080 27588
rect 24820 27548 24826 27560
rect 28074 27548 28080 27560
rect 28132 27548 28138 27600
rect 28166 27548 28172 27600
rect 28224 27588 28230 27600
rect 28308 27588 28336 27619
rect 28442 27616 28448 27668
rect 28500 27656 28506 27668
rect 31938 27656 31944 27668
rect 28500 27628 31944 27656
rect 28500 27616 28506 27628
rect 31938 27616 31944 27628
rect 31996 27616 32002 27668
rect 28224 27560 28336 27588
rect 28224 27548 28230 27560
rect 28534 27548 28540 27600
rect 28592 27588 28598 27600
rect 28718 27588 28724 27600
rect 28592 27560 28724 27588
rect 28592 27548 28598 27560
rect 28718 27548 28724 27560
rect 28776 27548 28782 27600
rect 31110 27588 31116 27600
rect 28966 27560 31116 27588
rect 23017 27523 23075 27529
rect 23017 27489 23029 27523
rect 23063 27489 23075 27523
rect 23017 27483 23075 27489
rect 25498 27480 25504 27532
rect 25556 27520 25562 27532
rect 25556 27492 26648 27520
rect 25556 27480 25562 27492
rect 20441 27455 20499 27461
rect 20441 27421 20453 27455
rect 20487 27421 20499 27455
rect 20441 27415 20499 27421
rect 21821 27455 21879 27461
rect 21821 27421 21833 27455
rect 21867 27421 21879 27455
rect 21821 27415 21879 27421
rect 20622 27384 20628 27396
rect 19444 27356 20628 27384
rect 19337 27347 19395 27353
rect 20622 27344 20628 27356
rect 20680 27344 20686 27396
rect 21082 27384 21088 27396
rect 21043 27356 21088 27384
rect 21082 27344 21088 27356
rect 21140 27344 21146 27396
rect 21726 27344 21732 27396
rect 21784 27384 21790 27396
rect 21836 27384 21864 27415
rect 21910 27412 21916 27464
rect 21968 27452 21974 27464
rect 22005 27455 22063 27461
rect 22005 27452 22017 27455
rect 21968 27424 22017 27452
rect 21968 27412 21974 27424
rect 22005 27421 22017 27424
rect 22051 27421 22063 27455
rect 23198 27452 23204 27464
rect 23159 27424 23204 27452
rect 22005 27415 22063 27421
rect 23198 27412 23204 27424
rect 23256 27412 23262 27464
rect 23934 27412 23940 27464
rect 23992 27452 23998 27464
rect 24394 27452 24400 27464
rect 23992 27424 24400 27452
rect 23992 27412 23998 27424
rect 24394 27412 24400 27424
rect 24452 27412 24458 27464
rect 24857 27455 24915 27461
rect 24857 27421 24869 27455
rect 24903 27452 24915 27455
rect 24946 27452 24952 27464
rect 24903 27424 24952 27452
rect 24903 27421 24915 27424
rect 24857 27415 24915 27421
rect 24946 27412 24952 27424
rect 25004 27452 25010 27464
rect 26510 27452 26516 27464
rect 25004 27424 26280 27452
rect 26471 27424 26516 27452
rect 25004 27412 25010 27424
rect 23014 27384 23020 27396
rect 21784 27356 23020 27384
rect 21784 27344 21790 27356
rect 23014 27344 23020 27356
rect 23072 27344 23078 27396
rect 23750 27344 23756 27396
rect 23808 27384 23814 27396
rect 25777 27387 25835 27393
rect 25777 27384 25789 27387
rect 23808 27356 25789 27384
rect 23808 27344 23814 27356
rect 25777 27353 25789 27356
rect 25823 27353 25835 27387
rect 26252 27384 26280 27424
rect 26510 27412 26516 27424
rect 26568 27412 26574 27464
rect 26620 27452 26648 27492
rect 26694 27480 26700 27532
rect 26752 27520 26758 27532
rect 28966 27520 28994 27560
rect 31110 27548 31116 27560
rect 31168 27548 31174 27600
rect 31846 27588 31852 27600
rect 31220 27560 31852 27588
rect 26752 27492 28994 27520
rect 29825 27523 29883 27529
rect 26752 27480 26758 27492
rect 29825 27489 29837 27523
rect 29871 27520 29883 27523
rect 30742 27520 30748 27532
rect 29871 27492 30748 27520
rect 29871 27489 29883 27492
rect 29825 27483 29883 27489
rect 30742 27480 30748 27492
rect 30800 27520 30806 27532
rect 31018 27520 31024 27532
rect 30800 27492 31024 27520
rect 30800 27480 30806 27492
rect 31018 27480 31024 27492
rect 31076 27480 31082 27532
rect 27157 27455 27215 27461
rect 27157 27452 27169 27455
rect 26620 27424 27169 27452
rect 27157 27421 27169 27424
rect 27203 27421 27215 27455
rect 27157 27415 27215 27421
rect 27341 27455 27399 27461
rect 27341 27421 27353 27455
rect 27387 27421 27399 27455
rect 27341 27415 27399 27421
rect 26252 27356 26740 27384
rect 25777 27347 25835 27353
rect 15473 27319 15531 27325
rect 15473 27285 15485 27319
rect 15519 27316 15531 27319
rect 16114 27316 16120 27328
rect 15519 27288 16120 27316
rect 15519 27285 15531 27288
rect 15473 27279 15531 27285
rect 16114 27276 16120 27288
rect 16172 27276 16178 27328
rect 17034 27276 17040 27328
rect 17092 27316 17098 27328
rect 17129 27319 17187 27325
rect 17129 27316 17141 27319
rect 17092 27288 17141 27316
rect 17092 27276 17098 27288
rect 17129 27285 17141 27288
rect 17175 27316 17187 27319
rect 18325 27319 18383 27325
rect 18325 27316 18337 27319
rect 17175 27288 18337 27316
rect 17175 27285 17187 27288
rect 17129 27279 17187 27285
rect 18325 27285 18337 27288
rect 18371 27285 18383 27319
rect 18325 27279 18383 27285
rect 18506 27276 18512 27328
rect 18564 27316 18570 27328
rect 20162 27316 20168 27328
rect 18564 27288 20168 27316
rect 18564 27276 18570 27288
rect 20162 27276 20168 27288
rect 20220 27316 20226 27328
rect 20349 27319 20407 27325
rect 20349 27316 20361 27319
rect 20220 27288 20361 27316
rect 20220 27276 20226 27288
rect 20349 27285 20361 27288
rect 20395 27285 20407 27319
rect 20349 27279 20407 27285
rect 20530 27276 20536 27328
rect 20588 27316 20594 27328
rect 22189 27319 22247 27325
rect 22189 27316 22201 27319
rect 20588 27288 22201 27316
rect 20588 27276 20594 27288
rect 22189 27285 22201 27288
rect 22235 27316 22247 27319
rect 22554 27316 22560 27328
rect 22235 27288 22560 27316
rect 22235 27285 22247 27288
rect 22189 27279 22247 27285
rect 22554 27276 22560 27288
rect 22612 27276 22618 27328
rect 23290 27276 23296 27328
rect 23348 27316 23354 27328
rect 23385 27319 23443 27325
rect 23385 27316 23397 27319
rect 23348 27288 23397 27316
rect 23348 27276 23354 27288
rect 23385 27285 23397 27288
rect 23431 27285 23443 27319
rect 23385 27279 23443 27285
rect 24210 27276 24216 27328
rect 24268 27316 24274 27328
rect 25133 27319 25191 27325
rect 25133 27316 25145 27319
rect 24268 27288 25145 27316
rect 24268 27276 24274 27288
rect 25133 27285 25145 27288
rect 25179 27316 25191 27319
rect 25682 27316 25688 27328
rect 25179 27288 25688 27316
rect 25179 27285 25191 27288
rect 25133 27279 25191 27285
rect 25682 27276 25688 27288
rect 25740 27276 25746 27328
rect 26602 27316 26608 27328
rect 26563 27288 26608 27316
rect 26602 27276 26608 27288
rect 26660 27276 26666 27328
rect 26712 27316 26740 27356
rect 26878 27344 26884 27396
rect 26936 27384 26942 27396
rect 27356 27384 27384 27415
rect 27430 27412 27436 27464
rect 27488 27452 27494 27464
rect 29362 27452 29368 27464
rect 27488 27424 29368 27452
rect 27488 27412 27494 27424
rect 29362 27412 29368 27424
rect 29420 27412 29426 27464
rect 29638 27452 29644 27464
rect 29599 27424 29644 27452
rect 29638 27412 29644 27424
rect 29696 27412 29702 27464
rect 29730 27412 29736 27464
rect 29788 27452 29794 27464
rect 30285 27455 30343 27461
rect 30285 27452 30297 27455
rect 29788 27424 30297 27452
rect 29788 27412 29794 27424
rect 30285 27421 30297 27424
rect 30331 27452 30343 27455
rect 30374 27452 30380 27464
rect 30331 27424 30380 27452
rect 30331 27421 30343 27424
rect 30285 27415 30343 27421
rect 30374 27412 30380 27424
rect 30432 27412 30438 27464
rect 30466 27412 30472 27464
rect 30524 27452 30530 27464
rect 30650 27452 30656 27464
rect 30524 27424 30656 27452
rect 30524 27412 30530 27424
rect 30650 27412 30656 27424
rect 30708 27412 30714 27464
rect 30834 27412 30840 27464
rect 30892 27452 30898 27464
rect 30929 27455 30987 27461
rect 30929 27452 30941 27455
rect 30892 27424 30941 27452
rect 30892 27412 30898 27424
rect 30929 27421 30941 27424
rect 30975 27421 30987 27455
rect 30929 27415 30987 27421
rect 26936 27356 27384 27384
rect 26936 27344 26942 27356
rect 27706 27344 27712 27396
rect 27764 27384 27770 27396
rect 27764 27356 27809 27384
rect 27764 27344 27770 27356
rect 27982 27344 27988 27396
rect 28040 27384 28046 27396
rect 28169 27387 28227 27393
rect 28169 27384 28181 27387
rect 28040 27356 28181 27384
rect 28040 27344 28046 27356
rect 28169 27353 28181 27356
rect 28215 27353 28227 27387
rect 31220 27384 31248 27560
rect 31846 27548 31852 27560
rect 31904 27548 31910 27600
rect 32306 27574 32312 27626
rect 32364 27574 32370 27626
rect 32398 27574 32404 27626
rect 32456 27574 32462 27626
rect 32490 27616 32496 27668
rect 32548 27656 32554 27668
rect 34514 27656 34520 27668
rect 32548 27628 34520 27656
rect 32548 27616 32554 27628
rect 34514 27616 34520 27628
rect 34572 27616 34578 27668
rect 34701 27591 34759 27597
rect 34701 27588 34713 27591
rect 31938 27520 31944 27532
rect 28169 27347 28227 27353
rect 28276 27356 31248 27384
rect 31404 27492 31944 27520
rect 28276 27316 28304 27356
rect 26712 27288 28304 27316
rect 28350 27276 28356 27328
rect 28408 27325 28414 27328
rect 28408 27319 28427 27325
rect 28415 27285 28427 27319
rect 28408 27279 28427 27285
rect 28408 27276 28414 27279
rect 28534 27276 28540 27328
rect 28592 27316 28598 27328
rect 30374 27316 30380 27328
rect 28592 27288 28637 27316
rect 30335 27288 30380 27316
rect 28592 27276 28598 27288
rect 30374 27276 30380 27288
rect 30432 27276 30438 27328
rect 30466 27276 30472 27328
rect 30524 27316 30530 27328
rect 31021 27319 31079 27325
rect 31021 27316 31033 27319
rect 30524 27288 31033 27316
rect 30524 27276 30530 27288
rect 31021 27285 31033 27288
rect 31067 27285 31079 27319
rect 31404 27316 31432 27492
rect 31938 27480 31944 27492
rect 31996 27480 32002 27532
rect 32030 27480 32036 27532
rect 32088 27520 32094 27532
rect 32125 27523 32183 27529
rect 32125 27520 32137 27523
rect 32088 27492 32137 27520
rect 32088 27480 32094 27492
rect 32125 27489 32137 27492
rect 32171 27489 32183 27523
rect 32125 27483 32183 27489
rect 31478 27412 31484 27464
rect 31536 27452 31542 27464
rect 31846 27452 31852 27464
rect 31536 27424 31852 27452
rect 31536 27412 31542 27424
rect 31846 27412 31852 27424
rect 31904 27412 31910 27464
rect 32324 27461 32352 27574
rect 32409 27529 32437 27574
rect 34164 27560 34713 27588
rect 34164 27529 34192 27560
rect 34701 27557 34713 27560
rect 34747 27557 34759 27591
rect 34701 27551 34759 27557
rect 36633 27591 36691 27597
rect 36633 27557 36645 27591
rect 36679 27588 36691 27591
rect 37458 27588 37464 27600
rect 36679 27560 37464 27588
rect 36679 27557 36691 27560
rect 36633 27551 36691 27557
rect 37458 27548 37464 27560
rect 37516 27548 37522 27600
rect 32401 27523 32459 27529
rect 32401 27489 32413 27523
rect 32447 27489 32459 27523
rect 32401 27483 32459 27489
rect 34149 27523 34207 27529
rect 34149 27489 34161 27523
rect 34195 27489 34207 27523
rect 34149 27483 34207 27489
rect 34422 27480 34428 27532
rect 34480 27520 34486 27532
rect 35529 27523 35587 27529
rect 34480 27492 34744 27520
rect 34480 27480 34486 27492
rect 32217 27455 32275 27461
rect 32217 27421 32229 27455
rect 32263 27421 32275 27455
rect 32217 27415 32275 27421
rect 32309 27455 32367 27461
rect 32309 27421 32321 27455
rect 32355 27421 32367 27455
rect 32309 27415 32367 27421
rect 31754 27344 31760 27396
rect 31812 27384 31818 27396
rect 32232 27384 32260 27415
rect 33226 27412 33232 27464
rect 33284 27452 33290 27464
rect 33630 27455 33688 27461
rect 33630 27452 33642 27455
rect 33284 27424 33642 27452
rect 33284 27412 33290 27424
rect 33630 27421 33642 27424
rect 33676 27421 33688 27455
rect 33630 27415 33688 27421
rect 34057 27455 34115 27461
rect 34057 27421 34069 27455
rect 34103 27452 34115 27455
rect 34606 27452 34612 27464
rect 34103 27424 34612 27452
rect 34103 27421 34115 27424
rect 34057 27415 34115 27421
rect 34606 27412 34612 27424
rect 34664 27412 34670 27464
rect 34716 27461 34744 27492
rect 35529 27489 35541 27523
rect 35575 27520 35587 27523
rect 35986 27520 35992 27532
rect 35575 27492 35992 27520
rect 35575 27489 35587 27492
rect 35529 27483 35587 27489
rect 35986 27480 35992 27492
rect 36044 27480 36050 27532
rect 36170 27520 36176 27532
rect 36131 27492 36176 27520
rect 36170 27480 36176 27492
rect 36228 27480 36234 27532
rect 36722 27480 36728 27532
rect 36780 27520 36786 27532
rect 36780 27492 37320 27520
rect 36780 27480 36786 27492
rect 34701 27455 34759 27461
rect 34701 27421 34713 27455
rect 34747 27421 34759 27455
rect 34701 27415 34759 27421
rect 35437 27455 35495 27461
rect 35437 27421 35449 27455
rect 35483 27421 35495 27455
rect 35618 27452 35624 27464
rect 35579 27424 35624 27452
rect 35437 27415 35495 27421
rect 35452 27384 35480 27415
rect 35618 27412 35624 27424
rect 35676 27412 35682 27464
rect 36265 27455 36323 27461
rect 36265 27421 36277 27455
rect 36311 27421 36323 27455
rect 36265 27415 36323 27421
rect 31812 27356 32260 27384
rect 33520 27356 35480 27384
rect 36280 27384 36308 27415
rect 36354 27412 36360 27464
rect 36412 27452 36418 27464
rect 37292 27461 37320 27492
rect 37093 27455 37151 27461
rect 37093 27452 37105 27455
rect 36412 27424 37105 27452
rect 36412 27412 36418 27424
rect 37093 27421 37105 27424
rect 37139 27421 37151 27455
rect 37093 27415 37151 27421
rect 37277 27455 37335 27461
rect 37277 27421 37289 27455
rect 37323 27421 37335 27455
rect 37734 27452 37740 27464
rect 37695 27424 37740 27452
rect 37277 27415 37335 27421
rect 37734 27412 37740 27424
rect 37792 27412 37798 27464
rect 37921 27455 37979 27461
rect 37921 27421 37933 27455
rect 37967 27452 37979 27455
rect 38102 27452 38108 27464
rect 37967 27424 38108 27452
rect 37967 27421 37979 27424
rect 37921 27415 37979 27421
rect 38102 27412 38108 27424
rect 38160 27412 38166 27464
rect 37185 27387 37243 27393
rect 37185 27384 37197 27387
rect 36280 27356 37197 27384
rect 31812 27344 31818 27356
rect 31478 27316 31484 27328
rect 31404 27288 31484 27316
rect 31021 27279 31079 27285
rect 31478 27276 31484 27288
rect 31536 27276 31542 27328
rect 31941 27319 31999 27325
rect 31941 27285 31953 27319
rect 31987 27316 31999 27319
rect 33410 27316 33416 27328
rect 31987 27288 33416 27316
rect 31987 27285 31999 27288
rect 31941 27279 31999 27285
rect 33410 27276 33416 27288
rect 33468 27276 33474 27328
rect 33520 27325 33548 27356
rect 37185 27353 37197 27356
rect 37231 27353 37243 27387
rect 37185 27347 37243 27353
rect 33505 27319 33563 27325
rect 33505 27285 33517 27319
rect 33551 27285 33563 27319
rect 33686 27316 33692 27328
rect 33647 27288 33692 27316
rect 33505 27279 33563 27285
rect 33686 27276 33692 27288
rect 33744 27276 33750 27328
rect 33778 27276 33784 27328
rect 33836 27316 33842 27328
rect 35066 27316 35072 27328
rect 33836 27288 35072 27316
rect 33836 27276 33842 27288
rect 35066 27276 35072 27288
rect 35124 27316 35130 27328
rect 36078 27316 36084 27328
rect 35124 27288 36084 27316
rect 35124 27276 35130 27288
rect 36078 27276 36084 27288
rect 36136 27276 36142 27328
rect 37274 27276 37280 27328
rect 37332 27316 37338 27328
rect 37829 27319 37887 27325
rect 37829 27316 37841 27319
rect 37332 27288 37841 27316
rect 37332 27276 37338 27288
rect 37829 27285 37841 27288
rect 37875 27285 37887 27319
rect 37829 27279 37887 27285
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 15381 27115 15439 27121
rect 15381 27081 15393 27115
rect 15427 27112 15439 27115
rect 15930 27112 15936 27124
rect 15427 27084 15936 27112
rect 15427 27081 15439 27084
rect 15381 27075 15439 27081
rect 15930 27072 15936 27084
rect 15988 27072 15994 27124
rect 20254 27112 20260 27124
rect 16776 27084 20260 27112
rect 16776 26988 16804 27084
rect 20254 27072 20260 27084
rect 20312 27072 20318 27124
rect 20346 27072 20352 27124
rect 20404 27112 20410 27124
rect 20404 27084 20449 27112
rect 20404 27072 20410 27084
rect 24854 27072 24860 27124
rect 24912 27112 24918 27124
rect 25041 27115 25099 27121
rect 25041 27112 25053 27115
rect 24912 27084 25053 27112
rect 24912 27072 24918 27084
rect 25041 27081 25053 27084
rect 25087 27081 25099 27115
rect 25041 27075 25099 27081
rect 25222 27072 25228 27124
rect 25280 27112 25286 27124
rect 25961 27115 26019 27121
rect 25961 27112 25973 27115
rect 25280 27084 25973 27112
rect 25280 27072 25286 27084
rect 25961 27081 25973 27084
rect 26007 27112 26019 27115
rect 26050 27112 26056 27124
rect 26007 27084 26056 27112
rect 26007 27081 26019 27084
rect 25961 27075 26019 27081
rect 26050 27072 26056 27084
rect 26108 27072 26114 27124
rect 28813 27115 28871 27121
rect 26160 27084 28580 27112
rect 18046 27044 18052 27056
rect 18007 27016 18052 27044
rect 18046 27004 18052 27016
rect 18104 27044 18110 27056
rect 19613 27047 19671 27053
rect 19613 27044 19625 27047
rect 18104 27016 19625 27044
rect 18104 27004 18110 27016
rect 19613 27013 19625 27016
rect 19659 27044 19671 27047
rect 20990 27044 20996 27056
rect 19659 27016 20996 27044
rect 19659 27013 19671 27016
rect 19613 27007 19671 27013
rect 20990 27004 20996 27016
rect 21048 27044 21054 27056
rect 21085 27047 21143 27053
rect 21085 27044 21097 27047
rect 21048 27016 21097 27044
rect 21048 27004 21054 27016
rect 21085 27013 21097 27016
rect 21131 27013 21143 27047
rect 21085 27007 21143 27013
rect 21269 27047 21327 27053
rect 21269 27013 21281 27047
rect 21315 27044 21327 27047
rect 22002 27044 22008 27056
rect 21315 27016 22008 27044
rect 21315 27013 21327 27016
rect 21269 27007 21327 27013
rect 22002 27004 22008 27016
rect 22060 27004 22066 27056
rect 23661 27047 23719 27053
rect 22204 27016 22692 27044
rect 14642 26976 14648 26988
rect 14603 26948 14648 26976
rect 14642 26936 14648 26948
rect 14700 26936 14706 26988
rect 15930 26976 15936 26988
rect 15891 26948 15936 26976
rect 15930 26936 15936 26948
rect 15988 26936 15994 26988
rect 16114 26976 16120 26988
rect 16075 26948 16120 26976
rect 16114 26936 16120 26948
rect 16172 26936 16178 26988
rect 16758 26976 16764 26988
rect 16671 26948 16764 26976
rect 16758 26936 16764 26948
rect 16816 26936 16822 26988
rect 17954 26936 17960 26988
rect 18012 26976 18018 26988
rect 19242 26976 19248 26988
rect 18012 26948 19248 26976
rect 18012 26936 18018 26948
rect 19242 26936 19248 26948
rect 19300 26976 19306 26988
rect 19429 26979 19487 26985
rect 19429 26976 19441 26979
rect 19300 26948 19441 26976
rect 19300 26936 19306 26948
rect 19429 26945 19441 26948
rect 19475 26945 19487 26979
rect 19429 26939 19487 26945
rect 19705 26979 19763 26985
rect 19705 26945 19717 26979
rect 19751 26945 19763 26979
rect 19705 26939 19763 26945
rect 14274 26868 14280 26920
rect 14332 26908 14338 26920
rect 14369 26911 14427 26917
rect 14369 26908 14381 26911
rect 14332 26880 14381 26908
rect 14332 26868 14338 26880
rect 14369 26877 14381 26880
rect 14415 26877 14427 26911
rect 14369 26871 14427 26877
rect 15286 26868 15292 26920
rect 15344 26908 15350 26920
rect 16853 26911 16911 26917
rect 16853 26908 16865 26911
rect 15344 26880 16865 26908
rect 15344 26868 15350 26880
rect 16853 26877 16865 26880
rect 16899 26908 16911 26911
rect 19518 26908 19524 26920
rect 16899 26880 19524 26908
rect 16899 26877 16911 26880
rect 16853 26871 16911 26877
rect 19518 26868 19524 26880
rect 19576 26868 19582 26920
rect 17681 26843 17739 26849
rect 17681 26809 17693 26843
rect 17727 26840 17739 26843
rect 18138 26840 18144 26852
rect 17727 26812 18144 26840
rect 17727 26809 17739 26812
rect 17681 26803 17739 26809
rect 18138 26800 18144 26812
rect 18196 26800 18202 26852
rect 18322 26800 18328 26852
rect 18380 26840 18386 26852
rect 19720 26840 19748 26939
rect 20070 26936 20076 26988
rect 20128 26976 20134 26988
rect 20165 26979 20223 26985
rect 20165 26976 20177 26979
rect 20128 26948 20177 26976
rect 20128 26936 20134 26948
rect 20165 26945 20177 26948
rect 20211 26945 20223 26979
rect 20165 26939 20223 26945
rect 20438 26936 20444 26988
rect 20496 26976 20502 26988
rect 20496 26948 20541 26976
rect 20496 26936 20502 26948
rect 20622 26936 20628 26988
rect 20680 26976 20686 26988
rect 22204 26976 22232 27016
rect 22370 26976 22376 26988
rect 20680 26948 22232 26976
rect 22331 26948 22376 26976
rect 20680 26936 20686 26948
rect 22370 26936 22376 26948
rect 22428 26936 22434 26988
rect 22664 26985 22692 27016
rect 23661 27013 23673 27047
rect 23707 27044 23719 27047
rect 24670 27044 24676 27056
rect 23707 27016 24676 27044
rect 23707 27013 23719 27016
rect 23661 27007 23719 27013
rect 24670 27004 24676 27016
rect 24728 27004 24734 27056
rect 25406 27004 25412 27056
rect 25464 27044 25470 27056
rect 26160 27044 26188 27084
rect 28442 27044 28448 27056
rect 25464 27016 26188 27044
rect 28403 27016 28448 27044
rect 25464 27004 25470 27016
rect 28442 27004 28448 27016
rect 28500 27004 28506 27056
rect 28552 27044 28580 27084
rect 28813 27081 28825 27115
rect 28859 27112 28871 27115
rect 33042 27112 33048 27124
rect 28859 27084 33048 27112
rect 28859 27081 28871 27084
rect 28813 27075 28871 27081
rect 33042 27072 33048 27084
rect 33100 27072 33106 27124
rect 33134 27072 33140 27124
rect 33192 27112 33198 27124
rect 33505 27115 33563 27121
rect 33505 27112 33517 27115
rect 33192 27084 33517 27112
rect 33192 27072 33198 27084
rect 33505 27081 33517 27084
rect 33551 27081 33563 27115
rect 33505 27075 33563 27081
rect 33781 27115 33839 27121
rect 33781 27081 33793 27115
rect 33827 27081 33839 27115
rect 33781 27075 33839 27081
rect 29730 27044 29736 27056
rect 28552 27016 29736 27044
rect 29730 27004 29736 27016
rect 29788 27004 29794 27056
rect 29917 27047 29975 27053
rect 29917 27013 29929 27047
rect 29963 27044 29975 27047
rect 30098 27044 30104 27056
rect 29963 27016 30104 27044
rect 29963 27013 29975 27016
rect 29917 27007 29975 27013
rect 30098 27004 30104 27016
rect 30156 27004 30162 27056
rect 32490 27044 32496 27056
rect 32451 27016 32496 27044
rect 32490 27004 32496 27016
rect 32548 27004 32554 27056
rect 33318 27004 33324 27056
rect 33376 27044 33382 27056
rect 33413 27047 33471 27053
rect 33413 27044 33425 27047
rect 33376 27016 33425 27044
rect 33376 27004 33382 27016
rect 33413 27013 33425 27016
rect 33459 27044 33471 27047
rect 33686 27044 33692 27056
rect 33459 27016 33692 27044
rect 33459 27013 33471 27016
rect 33413 27007 33471 27013
rect 33686 27004 33692 27016
rect 33744 27004 33750 27056
rect 33796 27044 33824 27075
rect 33870 27072 33876 27124
rect 33928 27112 33934 27124
rect 36541 27115 36599 27121
rect 36541 27112 36553 27115
rect 33928 27084 36553 27112
rect 33928 27072 33934 27084
rect 36541 27081 36553 27084
rect 36587 27081 36599 27115
rect 36541 27075 36599 27081
rect 35618 27044 35624 27056
rect 33796 27016 35624 27044
rect 22649 26979 22707 26985
rect 22649 26945 22661 26979
rect 22695 26976 22707 26979
rect 23477 26979 23535 26985
rect 23477 26976 23489 26979
rect 22695 26948 23489 26976
rect 22695 26945 22707 26948
rect 22649 26939 22707 26945
rect 23477 26945 23489 26948
rect 23523 26945 23535 26979
rect 23477 26939 23535 26945
rect 23566 26936 23572 26988
rect 23624 26976 23630 26988
rect 23750 26976 23756 26988
rect 23624 26948 23756 26976
rect 23624 26936 23630 26948
rect 23750 26936 23756 26948
rect 23808 26976 23814 26988
rect 24121 26979 24179 26985
rect 24121 26976 24133 26979
rect 23808 26948 24133 26976
rect 23808 26936 23814 26948
rect 24121 26945 24133 26948
rect 24167 26945 24179 26979
rect 24121 26939 24179 26945
rect 24213 26979 24271 26985
rect 24213 26945 24225 26979
rect 24259 26976 24271 26979
rect 24578 26976 24584 26988
rect 24259 26948 24584 26976
rect 24259 26945 24271 26948
rect 24213 26939 24271 26945
rect 24578 26936 24584 26948
rect 24636 26936 24642 26988
rect 24946 26976 24952 26988
rect 24907 26948 24952 26976
rect 24946 26936 24952 26948
rect 25004 26936 25010 26988
rect 25133 26979 25191 26985
rect 25133 26945 25145 26979
rect 25179 26976 25191 26979
rect 25314 26976 25320 26988
rect 25179 26948 25320 26976
rect 25179 26945 25191 26948
rect 25133 26939 25191 26945
rect 25314 26936 25320 26948
rect 25372 26936 25378 26988
rect 25498 26936 25504 26988
rect 25556 26976 25562 26988
rect 25593 26979 25651 26985
rect 25593 26976 25605 26979
rect 25556 26948 25605 26976
rect 25556 26936 25562 26948
rect 25593 26945 25605 26948
rect 25639 26945 25651 26979
rect 25593 26939 25651 26945
rect 25774 26936 25780 26988
rect 25832 26976 25838 26988
rect 25832 26948 25877 26976
rect 25832 26936 25838 26948
rect 27522 26936 27528 26988
rect 27580 26976 27586 26988
rect 28074 26976 28080 26988
rect 27580 26948 28080 26976
rect 27580 26936 27586 26948
rect 28074 26936 28080 26948
rect 28132 26976 28138 26988
rect 28261 26979 28319 26985
rect 28261 26976 28273 26979
rect 28132 26948 28273 26976
rect 28132 26936 28138 26948
rect 28261 26945 28273 26948
rect 28307 26945 28319 26979
rect 28261 26939 28319 26945
rect 28537 26979 28595 26985
rect 28537 26945 28549 26979
rect 28583 26945 28595 26979
rect 28537 26939 28595 26945
rect 28675 26979 28733 26985
rect 28675 26945 28687 26979
rect 28721 26976 28733 26979
rect 29638 26976 29644 26988
rect 28721 26948 28856 26976
rect 29599 26948 29644 26976
rect 28721 26945 28733 26948
rect 28675 26939 28733 26945
rect 20254 26868 20260 26920
rect 20312 26908 20318 26920
rect 22738 26908 22744 26920
rect 20312 26880 22744 26908
rect 20312 26868 20318 26880
rect 22738 26868 22744 26880
rect 22796 26868 22802 26920
rect 22925 26911 22983 26917
rect 22925 26877 22937 26911
rect 22971 26908 22983 26911
rect 23014 26908 23020 26920
rect 22971 26880 23020 26908
rect 22971 26877 22983 26880
rect 22925 26871 22983 26877
rect 23014 26868 23020 26880
rect 23072 26908 23078 26920
rect 25682 26908 25688 26920
rect 23072 26880 25688 26908
rect 23072 26868 23078 26880
rect 25682 26868 25688 26880
rect 25740 26868 25746 26920
rect 18380 26812 19748 26840
rect 18380 26800 18386 26812
rect 19978 26800 19984 26852
rect 20036 26840 20042 26852
rect 20165 26843 20223 26849
rect 20165 26840 20177 26843
rect 20036 26812 20177 26840
rect 20036 26800 20042 26812
rect 20165 26809 20177 26812
rect 20211 26809 20223 26843
rect 20165 26803 20223 26809
rect 25406 26800 25412 26852
rect 25464 26840 25470 26852
rect 25792 26840 25820 26936
rect 26970 26908 26976 26920
rect 26931 26880 26976 26908
rect 26970 26868 26976 26880
rect 27028 26868 27034 26920
rect 27249 26911 27307 26917
rect 27249 26877 27261 26911
rect 27295 26877 27307 26911
rect 27249 26871 27307 26877
rect 25464 26812 25820 26840
rect 27264 26840 27292 26871
rect 27430 26868 27436 26920
rect 27488 26908 27494 26920
rect 28350 26908 28356 26920
rect 27488 26880 28356 26908
rect 27488 26868 27494 26880
rect 28350 26868 28356 26880
rect 28408 26868 28414 26920
rect 28552 26840 28580 26939
rect 28828 26920 28856 26948
rect 29638 26936 29644 26948
rect 29696 26936 29702 26988
rect 29825 26979 29883 26985
rect 29825 26945 29837 26979
rect 29871 26945 29883 26979
rect 30006 26976 30012 26988
rect 29967 26948 30012 26976
rect 29825 26939 29883 26945
rect 28810 26868 28816 26920
rect 28868 26868 28874 26920
rect 28994 26868 29000 26920
rect 29052 26908 29058 26920
rect 29454 26908 29460 26920
rect 29052 26880 29460 26908
rect 29052 26868 29058 26880
rect 29454 26868 29460 26880
rect 29512 26908 29518 26920
rect 29840 26908 29868 26939
rect 30006 26936 30012 26948
rect 30064 26936 30070 26988
rect 30558 26936 30564 26988
rect 30616 26976 30622 26988
rect 30616 26948 30788 26976
rect 30616 26936 30622 26948
rect 30650 26908 30656 26920
rect 29512 26880 29868 26908
rect 30611 26880 30656 26908
rect 29512 26868 29518 26880
rect 30650 26868 30656 26880
rect 30708 26868 30714 26920
rect 30760 26908 30788 26948
rect 30834 26936 30840 26988
rect 30892 26976 30898 26988
rect 31138 26979 31196 26985
rect 31138 26976 31150 26979
rect 30892 26948 31150 26976
rect 30892 26936 30898 26948
rect 31138 26945 31150 26948
rect 31184 26945 31196 26979
rect 32214 26976 32220 26988
rect 31138 26939 31196 26945
rect 31312 26948 32220 26976
rect 30929 26911 30987 26917
rect 30929 26908 30941 26911
rect 30760 26880 30941 26908
rect 30929 26877 30941 26880
rect 30975 26877 30987 26911
rect 30929 26871 30987 26877
rect 31021 26911 31079 26917
rect 31021 26877 31033 26911
rect 31067 26908 31079 26911
rect 31312 26908 31340 26948
rect 32214 26936 32220 26948
rect 32272 26936 32278 26988
rect 32309 26979 32367 26985
rect 32309 26945 32321 26979
rect 32355 26945 32367 26979
rect 32309 26939 32367 26945
rect 31067 26880 31340 26908
rect 31067 26877 31079 26880
rect 31021 26871 31079 26877
rect 31386 26868 31392 26920
rect 31444 26908 31450 26920
rect 31570 26908 31576 26920
rect 31444 26880 31576 26908
rect 31444 26868 31450 26880
rect 31570 26868 31576 26880
rect 31628 26868 31634 26920
rect 31754 26868 31760 26920
rect 31812 26908 31818 26920
rect 32325 26908 32353 26939
rect 32398 26936 32404 26988
rect 32456 26976 32462 26988
rect 32677 26979 32735 26985
rect 32456 26948 32501 26976
rect 32456 26936 32462 26948
rect 32677 26945 32689 26979
rect 32723 26976 32735 26979
rect 33137 26979 33195 26985
rect 33137 26976 33149 26979
rect 32723 26948 33149 26976
rect 32723 26945 32735 26948
rect 32677 26939 32735 26945
rect 33137 26945 33149 26948
rect 33183 26976 33195 26979
rect 34606 26976 34612 26988
rect 33183 26948 34612 26976
rect 33183 26945 33195 26948
rect 33137 26939 33195 26945
rect 34606 26936 34612 26948
rect 34664 26936 34670 26988
rect 34716 26985 34744 27016
rect 35618 27004 35624 27016
rect 35676 27004 35682 27056
rect 34701 26979 34759 26985
rect 34701 26945 34713 26979
rect 34747 26945 34759 26979
rect 34701 26939 34759 26945
rect 34793 26979 34851 26985
rect 34793 26945 34805 26979
rect 34839 26945 34851 26979
rect 34793 26939 34851 26945
rect 34977 26979 35035 26985
rect 34977 26945 34989 26979
rect 35023 26976 35035 26979
rect 35066 26976 35072 26988
rect 35023 26948 35072 26976
rect 35023 26945 35035 26948
rect 34977 26939 35035 26945
rect 33502 26908 33508 26920
rect 31812 26880 33508 26908
rect 31812 26868 31818 26880
rect 33502 26868 33508 26880
rect 33560 26868 33566 26920
rect 33622 26911 33680 26917
rect 33622 26877 33634 26911
rect 33668 26908 33680 26911
rect 34422 26908 34428 26920
rect 33668 26880 34428 26908
rect 33668 26877 33680 26880
rect 33622 26871 33680 26877
rect 31846 26840 31852 26852
rect 27264 26812 31852 26840
rect 25464 26800 25470 26812
rect 31846 26800 31852 26812
rect 31904 26840 31910 26852
rect 32125 26843 32183 26849
rect 32125 26840 32137 26843
rect 31904 26812 32137 26840
rect 31904 26800 31910 26812
rect 32125 26809 32137 26812
rect 32171 26809 32183 26843
rect 32125 26803 32183 26809
rect 33042 26800 33048 26852
rect 33100 26840 33106 26852
rect 33637 26840 33665 26871
rect 34422 26868 34428 26880
rect 34480 26868 34486 26920
rect 34514 26840 34520 26852
rect 33100 26812 33665 26840
rect 34256 26812 34520 26840
rect 33100 26800 33106 26812
rect 15933 26775 15991 26781
rect 15933 26741 15945 26775
rect 15979 26772 15991 26775
rect 16666 26772 16672 26784
rect 15979 26744 16672 26772
rect 15979 26741 15991 26744
rect 15933 26735 15991 26741
rect 16666 26732 16672 26744
rect 16724 26732 16730 26784
rect 16850 26772 16856 26784
rect 16811 26744 16856 26772
rect 16850 26732 16856 26744
rect 16908 26732 16914 26784
rect 17129 26775 17187 26781
rect 17129 26741 17141 26775
rect 17175 26772 17187 26775
rect 17586 26772 17592 26784
rect 17175 26744 17592 26772
rect 17175 26741 17187 26744
rect 17129 26735 17187 26741
rect 17586 26732 17592 26744
rect 17644 26772 17650 26784
rect 17770 26772 17776 26784
rect 17644 26744 17776 26772
rect 17644 26732 17650 26744
rect 17770 26732 17776 26744
rect 17828 26732 17834 26784
rect 17954 26732 17960 26784
rect 18012 26772 18018 26784
rect 18049 26775 18107 26781
rect 18049 26772 18061 26775
rect 18012 26744 18061 26772
rect 18012 26732 18018 26744
rect 18049 26741 18061 26744
rect 18095 26741 18107 26775
rect 18230 26772 18236 26784
rect 18191 26744 18236 26772
rect 18049 26735 18107 26741
rect 18230 26732 18236 26744
rect 18288 26732 18294 26784
rect 19245 26775 19303 26781
rect 19245 26741 19257 26775
rect 19291 26772 19303 26775
rect 19886 26772 19892 26784
rect 19291 26744 19892 26772
rect 19291 26741 19303 26744
rect 19245 26735 19303 26741
rect 19886 26732 19892 26744
rect 19944 26732 19950 26784
rect 24302 26732 24308 26784
rect 24360 26772 24366 26784
rect 27522 26772 27528 26784
rect 24360 26744 27528 26772
rect 24360 26732 24366 26744
rect 27522 26732 27528 26744
rect 27580 26732 27586 26784
rect 28442 26732 28448 26784
rect 28500 26772 28506 26784
rect 29086 26772 29092 26784
rect 28500 26744 29092 26772
rect 28500 26732 28506 26744
rect 29086 26732 29092 26744
rect 29144 26732 29150 26784
rect 30193 26775 30251 26781
rect 30193 26741 30205 26775
rect 30239 26772 30251 26775
rect 30558 26772 30564 26784
rect 30239 26744 30564 26772
rect 30239 26741 30251 26744
rect 30193 26735 30251 26741
rect 30558 26732 30564 26744
rect 30616 26732 30622 26784
rect 31297 26775 31355 26781
rect 31297 26741 31309 26775
rect 31343 26772 31355 26775
rect 31478 26772 31484 26784
rect 31343 26744 31484 26772
rect 31343 26741 31355 26744
rect 31297 26735 31355 26741
rect 31478 26732 31484 26744
rect 31536 26732 31542 26784
rect 33226 26732 33232 26784
rect 33284 26772 33290 26784
rect 34256 26772 34284 26812
rect 34514 26800 34520 26812
rect 34572 26840 34578 26852
rect 34808 26840 34836 26939
rect 35066 26936 35072 26948
rect 35124 26936 35130 26988
rect 35710 26936 35716 26988
rect 35768 26976 35774 26988
rect 35768 26948 35813 26976
rect 35768 26936 35774 26948
rect 35894 26936 35900 26988
rect 35952 26976 35958 26988
rect 36446 26976 36452 26988
rect 35952 26948 35997 26976
rect 36407 26948 36452 26976
rect 35952 26936 35958 26948
rect 36446 26936 36452 26948
rect 36504 26936 36510 26988
rect 36538 26936 36544 26988
rect 36596 26976 36602 26988
rect 36633 26979 36691 26985
rect 36633 26976 36645 26979
rect 36596 26948 36645 26976
rect 36596 26936 36602 26948
rect 36633 26945 36645 26948
rect 36679 26945 36691 26979
rect 36633 26939 36691 26945
rect 37182 26936 37188 26988
rect 37240 26976 37246 26988
rect 37461 26979 37519 26985
rect 37461 26976 37473 26979
rect 37240 26948 37473 26976
rect 37240 26936 37246 26948
rect 37461 26945 37473 26948
rect 37507 26945 37519 26979
rect 37461 26939 37519 26945
rect 35618 26908 35624 26920
rect 35579 26880 35624 26908
rect 35618 26868 35624 26880
rect 35676 26868 35682 26920
rect 35805 26911 35863 26917
rect 35805 26877 35817 26911
rect 35851 26877 35863 26911
rect 37366 26908 37372 26920
rect 37327 26880 37372 26908
rect 35805 26871 35863 26877
rect 34572 26812 34836 26840
rect 35820 26840 35848 26871
rect 37366 26868 37372 26880
rect 37424 26868 37430 26920
rect 36722 26840 36728 26852
rect 35820 26812 36728 26840
rect 34572 26800 34578 26812
rect 36722 26800 36728 26812
rect 36780 26800 36786 26852
rect 33284 26744 34284 26772
rect 34333 26775 34391 26781
rect 33284 26732 33290 26744
rect 34333 26741 34345 26775
rect 34379 26772 34391 26775
rect 35342 26772 35348 26784
rect 34379 26744 35348 26772
rect 34379 26741 34391 26744
rect 34333 26735 34391 26741
rect 35342 26732 35348 26744
rect 35400 26732 35406 26784
rect 35437 26775 35495 26781
rect 35437 26741 35449 26775
rect 35483 26772 35495 26775
rect 36446 26772 36452 26784
rect 35483 26744 36452 26772
rect 35483 26741 35495 26744
rect 35437 26735 35495 26741
rect 36446 26732 36452 26744
rect 36504 26732 36510 26784
rect 37734 26772 37740 26784
rect 37695 26744 37740 26772
rect 37734 26732 37740 26744
rect 37792 26732 37798 26784
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 14274 26568 14280 26580
rect 14187 26540 14280 26568
rect 14200 26441 14228 26540
rect 14274 26528 14280 26540
rect 14332 26568 14338 26580
rect 15470 26568 15476 26580
rect 14332 26540 15476 26568
rect 14332 26528 14338 26540
rect 15470 26528 15476 26540
rect 15528 26528 15534 26580
rect 16758 26568 16764 26580
rect 16719 26540 16764 26568
rect 16758 26528 16764 26540
rect 16816 26528 16822 26580
rect 17770 26568 17776 26580
rect 17731 26540 17776 26568
rect 17770 26528 17776 26540
rect 17828 26528 17834 26580
rect 21910 26568 21916 26580
rect 18248 26540 21916 26568
rect 18248 26500 18276 26540
rect 17696 26472 18276 26500
rect 18325 26503 18383 26509
rect 14185 26435 14243 26441
rect 14185 26401 14197 26435
rect 14231 26401 14243 26435
rect 14185 26395 14243 26401
rect 14366 26324 14372 26376
rect 14424 26364 14430 26376
rect 14461 26367 14519 26373
rect 14461 26364 14473 26367
rect 14424 26336 14473 26364
rect 14424 26324 14430 26336
rect 14461 26333 14473 26336
rect 14507 26333 14519 26367
rect 15286 26364 15292 26376
rect 15247 26336 15292 26364
rect 14461 26327 14519 26333
rect 15286 26324 15292 26336
rect 15344 26324 15350 26376
rect 15470 26324 15476 26376
rect 15528 26364 15534 26376
rect 15749 26367 15807 26373
rect 15749 26364 15761 26367
rect 15528 26336 15761 26364
rect 15528 26324 15534 26336
rect 15749 26333 15761 26336
rect 15795 26333 15807 26367
rect 15749 26327 15807 26333
rect 16025 26367 16083 26373
rect 16025 26333 16037 26367
rect 16071 26333 16083 26367
rect 16025 26327 16083 26333
rect 13998 26256 14004 26308
rect 14056 26296 14062 26308
rect 16040 26296 16068 26327
rect 16666 26324 16672 26376
rect 16724 26364 16730 26376
rect 17696 26373 17724 26472
rect 18325 26469 18337 26503
rect 18371 26469 18383 26503
rect 18325 26463 18383 26469
rect 18049 26435 18107 26441
rect 18049 26401 18061 26435
rect 18095 26432 18107 26435
rect 18230 26432 18236 26444
rect 18095 26404 18236 26432
rect 18095 26401 18107 26404
rect 18049 26395 18107 26401
rect 18230 26392 18236 26404
rect 18288 26392 18294 26444
rect 18340 26432 18368 26463
rect 19334 26460 19340 26512
rect 19392 26500 19398 26512
rect 19705 26503 19763 26509
rect 19705 26500 19717 26503
rect 19392 26472 19717 26500
rect 19392 26460 19398 26472
rect 19705 26469 19717 26472
rect 19751 26469 19763 26503
rect 19705 26463 19763 26469
rect 21266 26432 21272 26444
rect 18340 26404 20208 26432
rect 20180 26376 20208 26404
rect 20732 26404 21272 26432
rect 20732 26376 20760 26404
rect 21266 26392 21272 26404
rect 21324 26392 21330 26444
rect 21450 26432 21456 26444
rect 21411 26404 21456 26432
rect 21450 26392 21456 26404
rect 21508 26392 21514 26444
rect 21836 26441 21864 26540
rect 21910 26528 21916 26540
rect 21968 26528 21974 26580
rect 24118 26528 24124 26580
rect 24176 26568 24182 26580
rect 25041 26571 25099 26577
rect 25041 26568 25053 26571
rect 24176 26540 25053 26568
rect 24176 26528 24182 26540
rect 25041 26537 25053 26540
rect 25087 26537 25099 26571
rect 25041 26531 25099 26537
rect 26697 26571 26755 26577
rect 26697 26537 26709 26571
rect 26743 26568 26755 26571
rect 26878 26568 26884 26580
rect 26743 26540 26884 26568
rect 26743 26537 26755 26540
rect 26697 26531 26755 26537
rect 26878 26528 26884 26540
rect 26936 26528 26942 26580
rect 27249 26571 27307 26577
rect 27249 26537 27261 26571
rect 27295 26568 27307 26571
rect 27706 26568 27712 26580
rect 27295 26540 27712 26568
rect 27295 26537 27307 26540
rect 27249 26531 27307 26537
rect 27706 26528 27712 26540
rect 27764 26528 27770 26580
rect 27798 26528 27804 26580
rect 27856 26528 27862 26580
rect 31754 26568 31760 26580
rect 28966 26540 31760 26568
rect 22462 26460 22468 26512
rect 22520 26500 22526 26512
rect 24136 26500 24164 26528
rect 22520 26472 24164 26500
rect 22520 26460 22526 26472
rect 25314 26460 25320 26512
rect 25372 26500 25378 26512
rect 26053 26503 26111 26509
rect 26053 26500 26065 26503
rect 25372 26472 26065 26500
rect 25372 26460 25378 26472
rect 26053 26469 26065 26472
rect 26099 26500 26111 26503
rect 26418 26500 26424 26512
rect 26099 26472 26424 26500
rect 26099 26469 26111 26472
rect 26053 26463 26111 26469
rect 26418 26460 26424 26472
rect 26476 26460 26482 26512
rect 26605 26503 26663 26509
rect 26605 26469 26617 26503
rect 26651 26500 26663 26503
rect 27816 26500 27844 26528
rect 26651 26472 27844 26500
rect 26651 26469 26663 26472
rect 26605 26463 26663 26469
rect 28166 26460 28172 26512
rect 28224 26500 28230 26512
rect 28537 26503 28595 26509
rect 28537 26500 28549 26503
rect 28224 26472 28549 26500
rect 28224 26460 28230 26472
rect 28537 26469 28549 26472
rect 28583 26500 28595 26503
rect 28966 26500 28994 26540
rect 31754 26528 31760 26540
rect 31812 26528 31818 26580
rect 33410 26528 33416 26580
rect 33468 26568 33474 26580
rect 35894 26568 35900 26580
rect 33468 26540 35756 26568
rect 35855 26540 35900 26568
rect 33468 26528 33474 26540
rect 28583 26472 28994 26500
rect 28583 26469 28595 26472
rect 28537 26463 28595 26469
rect 30650 26460 30656 26512
rect 30708 26500 30714 26512
rect 31570 26500 31576 26512
rect 30708 26472 31576 26500
rect 30708 26460 30714 26472
rect 31570 26460 31576 26472
rect 31628 26460 31634 26512
rect 33045 26503 33103 26509
rect 31680 26472 32996 26500
rect 21821 26435 21879 26441
rect 21821 26401 21833 26435
rect 21867 26401 21879 26435
rect 21821 26395 21879 26401
rect 23293 26435 23351 26441
rect 23293 26401 23305 26435
rect 23339 26432 23351 26435
rect 24210 26432 24216 26444
rect 23339 26404 24216 26432
rect 23339 26401 23351 26404
rect 23293 26395 23351 26401
rect 24210 26392 24216 26404
rect 24268 26392 24274 26444
rect 26789 26435 26847 26441
rect 25884 26404 26648 26432
rect 17681 26367 17739 26373
rect 17681 26364 17693 26367
rect 16724 26336 17693 26364
rect 16724 26324 16730 26336
rect 17681 26333 17693 26336
rect 17727 26333 17739 26367
rect 17681 26327 17739 26333
rect 18141 26367 18199 26373
rect 18141 26333 18153 26367
rect 18187 26333 18199 26367
rect 19886 26364 19892 26376
rect 19847 26336 19892 26364
rect 18141 26327 18199 26333
rect 14056 26268 16068 26296
rect 14056 26256 14062 26268
rect 16114 26256 16120 26308
rect 16172 26296 16178 26308
rect 18156 26296 18184 26327
rect 19886 26324 19892 26336
rect 19944 26324 19950 26376
rect 19981 26367 20039 26373
rect 19981 26333 19993 26367
rect 20027 26333 20039 26367
rect 20162 26364 20168 26376
rect 20075 26336 20168 26364
rect 19981 26327 20039 26333
rect 19996 26296 20024 26327
rect 20162 26324 20168 26336
rect 20220 26324 20226 26376
rect 20257 26367 20315 26373
rect 20257 26333 20269 26367
rect 20303 26364 20315 26367
rect 20714 26364 20720 26376
rect 20303 26336 20720 26364
rect 20303 26333 20315 26336
rect 20257 26327 20315 26333
rect 20714 26324 20720 26336
rect 20772 26324 20778 26376
rect 20990 26324 20996 26376
rect 21048 26364 21054 26376
rect 21545 26367 21603 26373
rect 21545 26364 21557 26367
rect 21048 26336 21557 26364
rect 21048 26324 21054 26336
rect 21545 26333 21557 26336
rect 21591 26333 21603 26367
rect 21910 26364 21916 26376
rect 21871 26336 21916 26364
rect 21545 26327 21603 26333
rect 21910 26324 21916 26336
rect 21968 26324 21974 26376
rect 23201 26367 23259 26373
rect 23201 26333 23213 26367
rect 23247 26364 23259 26367
rect 23382 26364 23388 26376
rect 23247 26336 23388 26364
rect 23247 26333 23259 26336
rect 23201 26327 23259 26333
rect 23382 26324 23388 26336
rect 23440 26364 23446 26376
rect 24302 26364 24308 26376
rect 23440 26336 24308 26364
rect 23440 26324 23446 26336
rect 24302 26324 24308 26336
rect 24360 26324 24366 26376
rect 25884 26373 25912 26404
rect 24949 26367 25007 26373
rect 24949 26333 24961 26367
rect 24995 26364 25007 26367
rect 25869 26367 25927 26373
rect 25869 26364 25881 26367
rect 24995 26336 25881 26364
rect 24995 26333 25007 26336
rect 24949 26327 25007 26333
rect 25869 26333 25881 26336
rect 25915 26333 25927 26367
rect 25869 26327 25927 26333
rect 26513 26367 26571 26373
rect 26513 26333 26525 26367
rect 26559 26333 26571 26367
rect 26620 26364 26648 26404
rect 26789 26401 26801 26435
rect 26835 26432 26847 26435
rect 27724 26432 27936 26440
rect 28994 26432 29000 26444
rect 26835 26412 29000 26432
rect 26835 26404 27752 26412
rect 27908 26404 29000 26412
rect 26835 26401 26847 26404
rect 26789 26395 26847 26401
rect 27062 26364 27068 26376
rect 26620 26336 27068 26364
rect 26513 26327 26571 26333
rect 20070 26296 20076 26308
rect 16172 26268 19932 26296
rect 19983 26268 20076 26296
rect 16172 26256 16178 26268
rect 19904 26228 19932 26268
rect 20070 26256 20076 26268
rect 20128 26296 20134 26308
rect 21269 26299 21327 26305
rect 21269 26296 21281 26299
rect 20128 26268 21281 26296
rect 20128 26256 20134 26268
rect 21269 26265 21281 26268
rect 21315 26265 21327 26299
rect 21269 26259 21327 26265
rect 23845 26299 23903 26305
rect 23845 26265 23857 26299
rect 23891 26296 23903 26299
rect 24394 26296 24400 26308
rect 23891 26268 24400 26296
rect 23891 26265 23903 26268
rect 23845 26259 23903 26265
rect 24394 26256 24400 26268
rect 24452 26256 24458 26308
rect 26528 26296 26556 26327
rect 27062 26324 27068 26336
rect 27120 26324 27126 26376
rect 27448 26373 27476 26404
rect 28994 26392 29000 26404
rect 29052 26392 29058 26444
rect 29178 26392 29184 26444
rect 29236 26432 29242 26444
rect 30745 26435 30803 26441
rect 30745 26432 30757 26435
rect 29236 26404 30757 26432
rect 29236 26392 29242 26404
rect 27433 26367 27491 26373
rect 27433 26333 27445 26367
rect 27479 26333 27491 26367
rect 27433 26327 27491 26333
rect 27522 26324 27528 26376
rect 27580 26364 27586 26376
rect 27709 26367 27767 26373
rect 27580 26336 27625 26364
rect 27580 26324 27586 26336
rect 27709 26333 27721 26367
rect 27755 26333 27767 26367
rect 27709 26327 27767 26333
rect 27724 26296 27752 26327
rect 27798 26324 27804 26376
rect 27856 26364 27862 26376
rect 28534 26364 28540 26376
rect 27856 26336 27901 26364
rect 28000 26336 28540 26364
rect 27856 26324 27862 26336
rect 28000 26296 28028 26336
rect 28534 26324 28540 26336
rect 28592 26324 28598 26376
rect 29564 26373 29592 26404
rect 30745 26401 30757 26404
rect 30791 26401 30803 26435
rect 31018 26432 31024 26444
rect 30745 26395 30803 26401
rect 30852 26404 31024 26432
rect 29549 26367 29607 26373
rect 29549 26333 29561 26367
rect 29595 26333 29607 26367
rect 29549 26327 29607 26333
rect 29733 26367 29791 26373
rect 29733 26333 29745 26367
rect 29779 26364 29791 26367
rect 30006 26364 30012 26376
rect 29779 26336 30012 26364
rect 29779 26333 29791 26336
rect 29733 26327 29791 26333
rect 30006 26324 30012 26336
rect 30064 26324 30070 26376
rect 30466 26364 30472 26376
rect 30427 26336 30472 26364
rect 30466 26324 30472 26336
rect 30524 26324 30530 26376
rect 30561 26367 30619 26373
rect 30561 26333 30573 26367
rect 30607 26364 30619 26367
rect 30650 26364 30656 26376
rect 30607 26336 30656 26364
rect 30607 26333 30619 26336
rect 30561 26327 30619 26333
rect 30650 26324 30656 26336
rect 30708 26324 30714 26376
rect 26528 26268 28028 26296
rect 28353 26299 28411 26305
rect 28353 26265 28365 26299
rect 28399 26296 28411 26299
rect 28810 26296 28816 26308
rect 28399 26268 28816 26296
rect 28399 26265 28411 26268
rect 28353 26259 28411 26265
rect 28810 26256 28816 26268
rect 28868 26256 28874 26308
rect 28994 26256 29000 26308
rect 29052 26296 29058 26308
rect 29641 26299 29699 26305
rect 29641 26296 29653 26299
rect 29052 26268 29653 26296
rect 29052 26256 29058 26268
rect 29641 26265 29653 26268
rect 29687 26265 29699 26299
rect 29641 26259 29699 26265
rect 30285 26299 30343 26305
rect 30285 26265 30297 26299
rect 30331 26296 30343 26299
rect 30374 26296 30380 26308
rect 30331 26268 30380 26296
rect 30331 26265 30343 26268
rect 30285 26259 30343 26265
rect 30374 26256 30380 26268
rect 30432 26256 30438 26308
rect 30760 26296 30788 26395
rect 30852 26373 30880 26404
rect 31018 26392 31024 26404
rect 31076 26392 31082 26444
rect 30837 26367 30895 26373
rect 30837 26333 30849 26367
rect 30883 26333 30895 26367
rect 30837 26327 30895 26333
rect 31680 26296 31708 26472
rect 31938 26392 31944 26444
rect 31996 26432 32002 26444
rect 32033 26435 32091 26441
rect 32033 26432 32045 26435
rect 31996 26404 32045 26432
rect 31996 26392 32002 26404
rect 32033 26401 32045 26404
rect 32079 26401 32091 26435
rect 32033 26395 32091 26401
rect 32582 26392 32588 26444
rect 32640 26432 32646 26444
rect 32968 26432 32996 26472
rect 33045 26469 33057 26503
rect 33091 26500 33103 26503
rect 34330 26500 34336 26512
rect 33091 26472 34336 26500
rect 33091 26469 33103 26472
rect 33045 26463 33103 26469
rect 34330 26460 34336 26472
rect 34388 26460 34394 26512
rect 34514 26460 34520 26512
rect 34572 26500 34578 26512
rect 34974 26500 34980 26512
rect 34572 26472 34980 26500
rect 34572 26460 34578 26472
rect 34974 26460 34980 26472
rect 35032 26460 35038 26512
rect 35728 26500 35756 26540
rect 35894 26528 35900 26540
rect 35952 26528 35958 26580
rect 36170 26568 36176 26580
rect 36131 26540 36176 26568
rect 36170 26528 36176 26540
rect 36228 26528 36234 26580
rect 37550 26500 37556 26512
rect 35728 26472 37556 26500
rect 37550 26460 37556 26472
rect 37608 26460 37614 26512
rect 33870 26432 33876 26444
rect 32640 26404 32904 26432
rect 32968 26404 33876 26432
rect 32640 26392 32646 26404
rect 32490 26364 32496 26376
rect 32451 26336 32496 26364
rect 32490 26324 32496 26336
rect 32548 26324 32554 26376
rect 32766 26364 32772 26376
rect 32600 26336 32772 26364
rect 31846 26296 31852 26308
rect 30760 26268 31708 26296
rect 31807 26268 31852 26296
rect 31846 26256 31852 26268
rect 31904 26296 31910 26308
rect 32600 26296 32628 26336
rect 32766 26324 32772 26336
rect 32824 26324 32830 26376
rect 32876 26373 32904 26404
rect 33870 26392 33876 26404
rect 33928 26392 33934 26444
rect 33965 26435 34023 26441
rect 33965 26401 33977 26435
rect 34011 26432 34023 26435
rect 34054 26432 34060 26444
rect 34011 26404 34060 26432
rect 34011 26401 34023 26404
rect 33965 26395 34023 26401
rect 34054 26392 34060 26404
rect 34112 26392 34118 26444
rect 34701 26435 34759 26441
rect 34701 26401 34713 26435
rect 34747 26432 34759 26435
rect 35618 26432 35624 26444
rect 34747 26404 35624 26432
rect 34747 26401 34759 26404
rect 34701 26395 34759 26401
rect 35618 26392 35624 26404
rect 35676 26432 35682 26444
rect 35676 26404 35756 26432
rect 35676 26392 35682 26404
rect 32861 26367 32919 26373
rect 32861 26333 32873 26367
rect 32907 26364 32919 26367
rect 33502 26364 33508 26376
rect 32907 26336 33508 26364
rect 32907 26333 32919 26336
rect 32861 26327 32919 26333
rect 33502 26324 33508 26336
rect 33560 26324 33566 26376
rect 34790 26324 34796 26376
rect 34848 26364 34854 26376
rect 34885 26367 34943 26373
rect 34885 26364 34897 26367
rect 34848 26336 34897 26364
rect 34848 26324 34854 26336
rect 34885 26333 34897 26336
rect 34931 26333 34943 26367
rect 34885 26327 34943 26333
rect 34974 26324 34980 26376
rect 35032 26364 35038 26376
rect 35161 26367 35219 26373
rect 35032 26336 35077 26364
rect 35032 26324 35038 26336
rect 35161 26333 35173 26367
rect 35207 26333 35219 26367
rect 35161 26327 35219 26333
rect 35253 26367 35311 26373
rect 35253 26333 35265 26367
rect 35299 26364 35311 26367
rect 35526 26364 35532 26376
rect 35299 26336 35532 26364
rect 35299 26333 35311 26336
rect 35253 26327 35311 26333
rect 31904 26268 32628 26296
rect 32677 26299 32735 26305
rect 31904 26256 31910 26268
rect 32677 26265 32689 26299
rect 32723 26296 32735 26299
rect 32723 26268 32812 26296
rect 32723 26265 32735 26268
rect 32677 26259 32735 26265
rect 21358 26228 21364 26240
rect 19904 26200 21364 26228
rect 21358 26188 21364 26200
rect 21416 26188 21422 26240
rect 21726 26228 21732 26240
rect 21687 26200 21732 26228
rect 21726 26188 21732 26200
rect 21784 26188 21790 26240
rect 23014 26188 23020 26240
rect 23072 26228 23078 26240
rect 27246 26228 27252 26240
rect 23072 26200 27252 26228
rect 23072 26188 23078 26200
rect 27246 26188 27252 26200
rect 27304 26188 27310 26240
rect 32784 26228 32812 26268
rect 33226 26256 33232 26308
rect 33284 26296 33290 26308
rect 33781 26299 33839 26305
rect 33781 26296 33793 26299
rect 33284 26268 33793 26296
rect 33284 26256 33290 26268
rect 33781 26265 33793 26268
rect 33827 26265 33839 26299
rect 33781 26259 33839 26265
rect 34606 26256 34612 26308
rect 34664 26296 34670 26308
rect 35176 26296 35204 26327
rect 35526 26324 35532 26336
rect 35584 26324 35590 26376
rect 35728 26373 35756 26404
rect 35713 26367 35771 26373
rect 35713 26333 35725 26367
rect 35759 26333 35771 26367
rect 35713 26327 35771 26333
rect 36446 26324 36452 26376
rect 36504 26364 36510 26376
rect 37277 26367 37335 26373
rect 37277 26364 37289 26367
rect 36504 26336 37289 26364
rect 36504 26324 36510 26336
rect 37277 26333 37289 26336
rect 37323 26333 37335 26367
rect 37734 26364 37740 26376
rect 37695 26336 37740 26364
rect 37277 26327 37335 26333
rect 37734 26324 37740 26336
rect 37792 26324 37798 26376
rect 34664 26268 35204 26296
rect 34664 26256 34670 26268
rect 37366 26256 37372 26308
rect 37424 26296 37430 26308
rect 38105 26299 38163 26305
rect 38105 26296 38117 26299
rect 37424 26268 38117 26296
rect 37424 26256 37430 26268
rect 38105 26265 38117 26268
rect 38151 26265 38163 26299
rect 38105 26259 38163 26265
rect 33042 26228 33048 26240
rect 32784 26200 33048 26228
rect 33042 26188 33048 26200
rect 33100 26188 33106 26240
rect 33502 26188 33508 26240
rect 33560 26228 33566 26240
rect 36538 26228 36544 26240
rect 33560 26200 36544 26228
rect 33560 26188 33566 26200
rect 36538 26188 36544 26200
rect 36596 26188 36602 26240
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 13173 26027 13231 26033
rect 13173 25993 13185 26027
rect 13219 26024 13231 26027
rect 14366 26024 14372 26036
rect 13219 25996 14372 26024
rect 13219 25993 13231 25996
rect 13173 25987 13231 25993
rect 14366 25984 14372 25996
rect 14424 25984 14430 26036
rect 14461 26027 14519 26033
rect 14461 25993 14473 26027
rect 14507 26024 14519 26027
rect 14642 26024 14648 26036
rect 14507 25996 14648 26024
rect 14507 25993 14519 25996
rect 14461 25987 14519 25993
rect 14642 25984 14648 25996
rect 14700 25984 14706 26036
rect 16114 26024 16120 26036
rect 16075 25996 16120 26024
rect 16114 25984 16120 25996
rect 16172 25984 16178 26036
rect 17681 26027 17739 26033
rect 17681 25993 17693 26027
rect 17727 26024 17739 26027
rect 17954 26024 17960 26036
rect 17727 25996 17960 26024
rect 17727 25993 17739 25996
rect 17681 25987 17739 25993
rect 17954 25984 17960 25996
rect 18012 25984 18018 26036
rect 18325 26027 18383 26033
rect 18325 25993 18337 26027
rect 18371 26024 18383 26027
rect 18506 26024 18512 26036
rect 18371 25996 18512 26024
rect 18371 25993 18383 25996
rect 18325 25987 18383 25993
rect 18506 25984 18512 25996
rect 18564 25984 18570 26036
rect 21450 25984 21456 26036
rect 21508 26024 21514 26036
rect 22557 26027 22615 26033
rect 22557 26024 22569 26027
rect 21508 25996 22569 26024
rect 21508 25984 21514 25996
rect 22557 25993 22569 25996
rect 22603 26024 22615 26027
rect 25590 26024 25596 26036
rect 22603 25996 25596 26024
rect 22603 25993 22615 25996
rect 22557 25987 22615 25993
rect 25590 25984 25596 25996
rect 25648 25984 25654 26036
rect 25866 25984 25872 26036
rect 25924 26024 25930 26036
rect 26602 26024 26608 26036
rect 25924 25996 26608 26024
rect 25924 25984 25930 25996
rect 26602 25984 26608 25996
rect 26660 25984 26666 26036
rect 28350 25984 28356 26036
rect 28408 26024 28414 26036
rect 30006 26024 30012 26036
rect 28408 25996 30012 26024
rect 28408 25984 28414 25996
rect 30006 25984 30012 25996
rect 30064 26024 30070 26036
rect 30561 26027 30619 26033
rect 30561 26024 30573 26027
rect 30064 25996 30573 26024
rect 30064 25984 30070 25996
rect 30561 25993 30573 25996
rect 30607 25993 30619 26027
rect 32030 26024 32036 26036
rect 30561 25987 30619 25993
rect 30668 25996 32036 26024
rect 15194 25956 15200 25968
rect 14016 25928 15200 25956
rect 13357 25891 13415 25897
rect 13357 25857 13369 25891
rect 13403 25888 13415 25891
rect 13906 25888 13912 25900
rect 13403 25860 13912 25888
rect 13403 25857 13415 25860
rect 13357 25851 13415 25857
rect 13906 25848 13912 25860
rect 13964 25848 13970 25900
rect 14016 25897 14044 25928
rect 15194 25916 15200 25928
rect 15252 25916 15258 25968
rect 18138 25916 18144 25968
rect 18196 25956 18202 25968
rect 18233 25959 18291 25965
rect 18233 25956 18245 25959
rect 18196 25928 18245 25956
rect 18196 25916 18202 25928
rect 18233 25925 18245 25928
rect 18279 25956 18291 25959
rect 18279 25928 18920 25956
rect 18279 25925 18291 25928
rect 18233 25919 18291 25925
rect 14001 25891 14059 25897
rect 14001 25857 14013 25891
rect 14047 25857 14059 25891
rect 14642 25888 14648 25900
rect 14603 25860 14648 25888
rect 14001 25851 14059 25857
rect 14642 25848 14648 25860
rect 14700 25848 14706 25900
rect 15378 25888 15384 25900
rect 15339 25860 15384 25888
rect 15378 25848 15384 25860
rect 15436 25848 15442 25900
rect 15746 25848 15752 25900
rect 15804 25888 15810 25900
rect 18892 25897 18920 25928
rect 19242 25916 19248 25968
rect 19300 25956 19306 25968
rect 24121 25959 24179 25965
rect 19300 25928 20760 25956
rect 19300 25916 19306 25928
rect 16945 25891 17003 25897
rect 16945 25888 16957 25891
rect 15804 25860 16957 25888
rect 15804 25848 15810 25860
rect 16945 25857 16957 25860
rect 16991 25857 17003 25891
rect 16945 25851 17003 25857
rect 18877 25891 18935 25897
rect 18877 25857 18889 25891
rect 18923 25857 18935 25891
rect 18877 25851 18935 25857
rect 19889 25891 19947 25897
rect 19889 25857 19901 25891
rect 19935 25888 19947 25891
rect 20070 25888 20076 25900
rect 19935 25860 20076 25888
rect 19935 25857 19947 25860
rect 19889 25851 19947 25857
rect 20070 25848 20076 25860
rect 20128 25848 20134 25900
rect 20162 25848 20168 25900
rect 20220 25888 20226 25900
rect 20732 25897 20760 25928
rect 24121 25925 24133 25959
rect 24167 25956 24179 25959
rect 25498 25956 25504 25968
rect 24167 25928 25504 25956
rect 24167 25925 24179 25928
rect 24121 25919 24179 25925
rect 25498 25916 25504 25928
rect 25556 25956 25562 25968
rect 27430 25956 27436 25968
rect 25556 25928 26372 25956
rect 27391 25928 27436 25956
rect 25556 25916 25562 25928
rect 20257 25891 20315 25897
rect 20257 25888 20269 25891
rect 20220 25860 20269 25888
rect 20220 25848 20226 25860
rect 20257 25857 20269 25860
rect 20303 25857 20315 25891
rect 20257 25851 20315 25857
rect 20717 25891 20775 25897
rect 20717 25857 20729 25891
rect 20763 25857 20775 25891
rect 20717 25851 20775 25857
rect 20901 25891 20959 25897
rect 20901 25857 20913 25891
rect 20947 25888 20959 25891
rect 21358 25888 21364 25900
rect 20947 25860 21364 25888
rect 20947 25857 20959 25860
rect 20901 25851 20959 25857
rect 21358 25848 21364 25860
rect 21416 25848 21422 25900
rect 22370 25888 22376 25900
rect 22331 25860 22376 25888
rect 22370 25848 22376 25860
rect 22428 25888 22434 25900
rect 23014 25888 23020 25900
rect 22428 25860 23020 25888
rect 22428 25848 22434 25860
rect 23014 25848 23020 25860
rect 23072 25888 23078 25900
rect 23109 25891 23167 25897
rect 23109 25888 23121 25891
rect 23072 25860 23121 25888
rect 23072 25848 23078 25860
rect 23109 25857 23121 25860
rect 23155 25857 23167 25891
rect 23109 25851 23167 25857
rect 23934 25848 23940 25900
rect 23992 25888 23998 25900
rect 24029 25891 24087 25897
rect 24029 25888 24041 25891
rect 23992 25860 24041 25888
rect 23992 25848 23998 25860
rect 24029 25857 24041 25860
rect 24075 25857 24087 25891
rect 24029 25851 24087 25857
rect 24213 25891 24271 25897
rect 24213 25857 24225 25891
rect 24259 25888 24271 25891
rect 24578 25888 24584 25900
rect 24259 25860 24584 25888
rect 24259 25857 24271 25860
rect 24213 25851 24271 25857
rect 15105 25823 15163 25829
rect 15105 25789 15117 25823
rect 15151 25789 15163 25823
rect 15105 25783 15163 25789
rect 13814 25752 13820 25764
rect 13775 25724 13820 25752
rect 13814 25712 13820 25724
rect 13872 25712 13878 25764
rect 15120 25684 15148 25783
rect 16390 25780 16396 25832
rect 16448 25820 16454 25832
rect 16669 25823 16727 25829
rect 16669 25820 16681 25823
rect 16448 25792 16681 25820
rect 16448 25780 16454 25792
rect 16669 25789 16681 25792
rect 16715 25789 16727 25823
rect 16669 25783 16727 25789
rect 19705 25823 19763 25829
rect 19705 25789 19717 25823
rect 19751 25820 19763 25823
rect 19978 25820 19984 25832
rect 19751 25792 19984 25820
rect 19751 25789 19763 25792
rect 19705 25783 19763 25789
rect 19978 25780 19984 25792
rect 20036 25780 20042 25832
rect 20809 25823 20867 25829
rect 20809 25789 20821 25823
rect 20855 25820 20867 25823
rect 21910 25820 21916 25832
rect 20855 25792 21916 25820
rect 20855 25789 20867 25792
rect 20809 25783 20867 25789
rect 21910 25780 21916 25792
rect 21968 25780 21974 25832
rect 22278 25780 22284 25832
rect 22336 25820 22342 25832
rect 24228 25820 24256 25851
rect 24578 25848 24584 25860
rect 24636 25848 24642 25900
rect 24857 25891 24915 25897
rect 24857 25857 24869 25891
rect 24903 25888 24915 25891
rect 24903 25860 25820 25888
rect 24903 25857 24915 25860
rect 24857 25851 24915 25857
rect 22336 25792 24256 25820
rect 22336 25780 22342 25792
rect 24394 25780 24400 25832
rect 24452 25820 24458 25832
rect 24949 25823 25007 25829
rect 24949 25820 24961 25823
rect 24452 25792 24961 25820
rect 24452 25780 24458 25792
rect 24949 25789 24961 25792
rect 24995 25789 25007 25823
rect 24949 25783 25007 25789
rect 25041 25823 25099 25829
rect 25041 25789 25053 25823
rect 25087 25789 25099 25823
rect 25041 25783 25099 25789
rect 25133 25823 25191 25829
rect 25133 25789 25145 25823
rect 25179 25820 25191 25823
rect 25222 25820 25228 25832
rect 25179 25792 25228 25820
rect 25179 25789 25191 25792
rect 25133 25783 25191 25789
rect 20165 25755 20223 25761
rect 20165 25721 20177 25755
rect 20211 25752 20223 25755
rect 20346 25752 20352 25764
rect 20211 25724 20352 25752
rect 20211 25721 20223 25724
rect 20165 25715 20223 25721
rect 20346 25712 20352 25724
rect 20404 25712 20410 25764
rect 23293 25755 23351 25761
rect 23293 25721 23305 25755
rect 23339 25752 23351 25755
rect 23382 25752 23388 25764
rect 23339 25724 23388 25752
rect 23339 25721 23351 25724
rect 23293 25715 23351 25721
rect 23382 25712 23388 25724
rect 23440 25712 23446 25764
rect 23842 25712 23848 25764
rect 23900 25752 23906 25764
rect 25056 25752 25084 25783
rect 25222 25780 25228 25792
rect 25280 25780 25286 25832
rect 25792 25820 25820 25860
rect 25866 25848 25872 25900
rect 25924 25888 25930 25900
rect 25924 25860 25969 25888
rect 25924 25848 25930 25860
rect 26050 25848 26056 25900
rect 26108 25888 26114 25900
rect 26344 25897 26372 25928
rect 27430 25916 27436 25928
rect 27488 25916 27494 25968
rect 27617 25959 27675 25965
rect 27617 25925 27629 25959
rect 27663 25956 27675 25959
rect 27982 25956 27988 25968
rect 27663 25928 27988 25956
rect 27663 25925 27675 25928
rect 27617 25919 27675 25925
rect 27982 25916 27988 25928
rect 28040 25956 28046 25968
rect 28902 25956 28908 25968
rect 28040 25928 28908 25956
rect 28040 25916 28046 25928
rect 28902 25916 28908 25928
rect 28960 25916 28966 25968
rect 29086 25916 29092 25968
rect 29144 25956 29150 25968
rect 29362 25956 29368 25968
rect 29144 25928 29368 25956
rect 29144 25916 29150 25928
rect 29362 25916 29368 25928
rect 29420 25916 29426 25968
rect 29581 25959 29639 25965
rect 29581 25925 29593 25959
rect 29627 25956 29639 25959
rect 29627 25928 30328 25956
rect 29627 25925 29639 25928
rect 29581 25919 29639 25925
rect 30300 25900 30328 25928
rect 26145 25891 26203 25897
rect 26145 25888 26157 25891
rect 26108 25860 26157 25888
rect 26108 25848 26114 25860
rect 26145 25857 26157 25860
rect 26191 25857 26203 25891
rect 26145 25851 26203 25857
rect 26329 25891 26387 25897
rect 26329 25857 26341 25891
rect 26375 25857 26387 25891
rect 26329 25851 26387 25857
rect 26510 25848 26516 25900
rect 26568 25888 26574 25900
rect 26786 25888 26792 25900
rect 26568 25860 26792 25888
rect 26568 25848 26574 25860
rect 26786 25848 26792 25860
rect 26844 25888 26850 25900
rect 27709 25891 27767 25897
rect 27709 25888 27721 25891
rect 26844 25860 27721 25888
rect 26844 25848 26850 25860
rect 27709 25857 27721 25860
rect 27755 25857 27767 25891
rect 27709 25851 27767 25857
rect 28537 25891 28595 25897
rect 28537 25857 28549 25891
rect 28583 25888 28595 25891
rect 29730 25888 29736 25900
rect 28583 25860 29736 25888
rect 28583 25857 28595 25860
rect 28537 25851 28595 25857
rect 29730 25848 29736 25860
rect 29788 25888 29794 25900
rect 30098 25888 30104 25900
rect 29788 25860 30104 25888
rect 29788 25848 29794 25860
rect 30098 25848 30104 25860
rect 30156 25848 30162 25900
rect 30282 25848 30288 25900
rect 30340 25888 30346 25900
rect 30668 25897 30696 25996
rect 32030 25984 32036 25996
rect 32088 25984 32094 26036
rect 32490 25984 32496 26036
rect 32548 26024 32554 26036
rect 33689 26027 33747 26033
rect 33689 26024 33701 26027
rect 32548 25996 33701 26024
rect 32548 25984 32554 25996
rect 33689 25993 33701 25996
rect 33735 25993 33747 26027
rect 33689 25987 33747 25993
rect 33778 25984 33784 26036
rect 33836 26024 33842 26036
rect 35345 26027 35403 26033
rect 35345 26024 35357 26027
rect 33836 25996 35357 26024
rect 33836 25984 33842 25996
rect 35345 25993 35357 25996
rect 35391 26024 35403 26027
rect 36722 26024 36728 26036
rect 35391 25996 36728 26024
rect 35391 25993 35403 25996
rect 35345 25987 35403 25993
rect 36722 25984 36728 25996
rect 36780 25984 36786 26036
rect 30926 25916 30932 25968
rect 30984 25956 30990 25968
rect 30984 25928 31754 25956
rect 30984 25916 30990 25928
rect 30377 25891 30435 25897
rect 30377 25888 30389 25891
rect 30340 25860 30389 25888
rect 30340 25848 30346 25860
rect 30377 25857 30389 25860
rect 30423 25857 30435 25891
rect 30377 25851 30435 25857
rect 30653 25891 30711 25897
rect 30653 25857 30665 25891
rect 30699 25857 30711 25891
rect 30653 25851 30711 25857
rect 30834 25848 30840 25900
rect 30892 25848 30898 25900
rect 31018 25848 31024 25900
rect 31076 25888 31082 25900
rect 31113 25891 31171 25897
rect 31113 25888 31125 25891
rect 31076 25860 31125 25888
rect 31076 25848 31082 25860
rect 31113 25857 31125 25860
rect 31159 25857 31171 25891
rect 31294 25888 31300 25900
rect 31255 25860 31300 25888
rect 31113 25851 31171 25857
rect 31294 25848 31300 25860
rect 31352 25848 31358 25900
rect 26234 25820 26240 25832
rect 25792 25792 26240 25820
rect 26234 25780 26240 25792
rect 26292 25780 26298 25832
rect 28626 25780 28632 25832
rect 28684 25820 28690 25832
rect 28721 25823 28779 25829
rect 28721 25820 28733 25823
rect 28684 25792 28733 25820
rect 28684 25780 28690 25792
rect 28721 25789 28733 25792
rect 28767 25789 28779 25823
rect 28721 25783 28779 25789
rect 28810 25780 28816 25832
rect 28868 25820 28874 25832
rect 30193 25823 30251 25829
rect 28868 25792 28913 25820
rect 28868 25780 28874 25792
rect 30193 25789 30205 25823
rect 30239 25820 30251 25823
rect 30852 25820 30880 25848
rect 30239 25792 30880 25820
rect 30239 25789 30251 25792
rect 30193 25783 30251 25789
rect 31386 25780 31392 25832
rect 31444 25780 31450 25832
rect 31726 25820 31754 25928
rect 31938 25916 31944 25968
rect 31996 25956 32002 25968
rect 32585 25959 32643 25965
rect 32585 25956 32597 25959
rect 31996 25928 32597 25956
rect 31996 25916 32002 25928
rect 32585 25925 32597 25928
rect 32631 25925 32643 25959
rect 32585 25919 32643 25925
rect 32766 25916 32772 25968
rect 32824 25956 32830 25968
rect 33321 25959 33379 25965
rect 33321 25956 33333 25959
rect 32824 25928 33333 25956
rect 32824 25916 32830 25928
rect 33321 25925 33333 25928
rect 33367 25925 33379 25959
rect 33502 25956 33508 25968
rect 33463 25928 33508 25956
rect 33321 25919 33379 25925
rect 33502 25916 33508 25928
rect 33560 25916 33566 25968
rect 35253 25959 35311 25965
rect 35253 25925 35265 25959
rect 35299 25956 35311 25959
rect 35710 25956 35716 25968
rect 35299 25928 35716 25956
rect 35299 25925 35311 25928
rect 35253 25919 35311 25925
rect 35710 25916 35716 25928
rect 35768 25956 35774 25968
rect 36081 25959 36139 25965
rect 36081 25956 36093 25959
rect 35768 25928 36093 25956
rect 35768 25916 35774 25928
rect 36081 25925 36093 25928
rect 36127 25925 36139 25959
rect 36081 25919 36139 25925
rect 32306 25888 32312 25900
rect 32267 25860 32312 25888
rect 32306 25848 32312 25860
rect 32364 25848 32370 25900
rect 32493 25891 32551 25897
rect 32493 25857 32505 25891
rect 32539 25857 32551 25891
rect 32493 25851 32551 25857
rect 32677 25891 32735 25897
rect 32677 25857 32689 25891
rect 32723 25888 32735 25891
rect 32950 25888 32956 25900
rect 32723 25860 32956 25888
rect 32723 25857 32735 25860
rect 32677 25851 32735 25857
rect 32508 25820 32536 25851
rect 32950 25848 32956 25860
rect 33008 25848 33014 25900
rect 33134 25848 33140 25900
rect 33192 25888 33198 25900
rect 33597 25891 33655 25897
rect 33597 25888 33609 25891
rect 33192 25860 33609 25888
rect 33192 25848 33198 25860
rect 33597 25857 33609 25860
rect 33643 25857 33655 25891
rect 34330 25888 34336 25900
rect 34291 25860 34336 25888
rect 33597 25851 33655 25857
rect 34330 25848 34336 25860
rect 34388 25848 34394 25900
rect 35897 25891 35955 25897
rect 35897 25857 35909 25891
rect 35943 25888 35955 25891
rect 35986 25888 35992 25900
rect 35943 25860 35992 25888
rect 35943 25857 35955 25860
rect 35897 25851 35955 25857
rect 35986 25848 35992 25860
rect 36044 25848 36050 25900
rect 36170 25888 36176 25900
rect 36131 25860 36176 25888
rect 36170 25848 36176 25860
rect 36228 25848 36234 25900
rect 37458 25888 37464 25900
rect 37419 25860 37464 25888
rect 37458 25848 37464 25860
rect 37516 25848 37522 25900
rect 37550 25820 37556 25832
rect 31726 25792 32536 25820
rect 37511 25792 37556 25820
rect 37550 25780 37556 25792
rect 37608 25780 37614 25832
rect 23900 25724 25084 25752
rect 23900 25712 23906 25724
rect 25866 25712 25872 25764
rect 25924 25752 25930 25764
rect 25961 25755 26019 25761
rect 25961 25752 25973 25755
rect 25924 25724 25973 25752
rect 25924 25712 25930 25724
rect 25961 25721 25973 25724
rect 26007 25721 26019 25755
rect 25961 25715 26019 25721
rect 26050 25712 26056 25764
rect 26108 25752 26114 25764
rect 27433 25755 27491 25761
rect 26108 25724 26153 25752
rect 26108 25712 26114 25724
rect 27433 25721 27445 25755
rect 27479 25752 27491 25755
rect 27798 25752 27804 25764
rect 27479 25724 27804 25752
rect 27479 25721 27491 25724
rect 27433 25715 27491 25721
rect 27798 25712 27804 25724
rect 27856 25712 27862 25764
rect 29733 25755 29791 25761
rect 29733 25721 29745 25755
rect 29779 25752 29791 25755
rect 30650 25752 30656 25764
rect 29779 25724 30656 25752
rect 29779 25721 29791 25724
rect 29733 25715 29791 25721
rect 30650 25712 30656 25724
rect 30708 25712 30714 25764
rect 31404 25752 31432 25780
rect 31662 25752 31668 25764
rect 31404 25724 31668 25752
rect 31662 25712 31668 25724
rect 31720 25712 31726 25764
rect 15470 25684 15476 25696
rect 15120 25656 15476 25684
rect 15470 25644 15476 25656
rect 15528 25644 15534 25696
rect 18322 25644 18328 25696
rect 18380 25684 18386 25696
rect 19058 25684 19064 25696
rect 18380 25656 19064 25684
rect 18380 25644 18386 25656
rect 19058 25644 19064 25656
rect 19116 25644 19122 25696
rect 23106 25644 23112 25696
rect 23164 25684 23170 25696
rect 23566 25684 23572 25696
rect 23164 25656 23572 25684
rect 23164 25644 23170 25656
rect 23566 25644 23572 25656
rect 23624 25644 23630 25696
rect 24673 25687 24731 25693
rect 24673 25653 24685 25687
rect 24719 25684 24731 25687
rect 25590 25684 25596 25696
rect 24719 25656 25596 25684
rect 24719 25653 24731 25656
rect 24673 25647 24731 25653
rect 25590 25644 25596 25656
rect 25648 25644 25654 25696
rect 25685 25687 25743 25693
rect 25685 25653 25697 25687
rect 25731 25684 25743 25687
rect 26418 25684 26424 25696
rect 25731 25656 26424 25684
rect 25731 25653 25743 25656
rect 25685 25647 25743 25653
rect 26418 25644 26424 25656
rect 26476 25644 26482 25696
rect 28353 25687 28411 25693
rect 28353 25653 28365 25687
rect 28399 25684 28411 25687
rect 28534 25684 28540 25696
rect 28399 25656 28540 25684
rect 28399 25653 28411 25656
rect 28353 25647 28411 25653
rect 28534 25644 28540 25656
rect 28592 25644 28598 25696
rect 29549 25687 29607 25693
rect 29549 25653 29561 25687
rect 29595 25684 29607 25687
rect 29914 25684 29920 25696
rect 29595 25656 29920 25684
rect 29595 25653 29607 25656
rect 29549 25647 29607 25653
rect 29914 25644 29920 25656
rect 29972 25644 29978 25696
rect 30282 25644 30288 25696
rect 30340 25684 30346 25696
rect 30742 25684 30748 25696
rect 30340 25656 30748 25684
rect 30340 25644 30346 25656
rect 30742 25644 30748 25656
rect 30800 25644 30806 25696
rect 31205 25687 31263 25693
rect 31205 25653 31217 25687
rect 31251 25684 31263 25687
rect 31386 25684 31392 25696
rect 31251 25656 31392 25684
rect 31251 25653 31263 25656
rect 31205 25647 31263 25653
rect 31386 25644 31392 25656
rect 31444 25644 31450 25696
rect 32490 25644 32496 25696
rect 32548 25684 32554 25696
rect 32861 25687 32919 25693
rect 32861 25684 32873 25687
rect 32548 25656 32873 25684
rect 32548 25644 32554 25656
rect 32861 25653 32873 25656
rect 32907 25653 32919 25687
rect 33870 25684 33876 25696
rect 33831 25656 33876 25684
rect 32861 25647 32919 25653
rect 33870 25644 33876 25656
rect 33928 25644 33934 25696
rect 34514 25684 34520 25696
rect 34475 25656 34520 25684
rect 34514 25644 34520 25656
rect 34572 25644 34578 25696
rect 35894 25684 35900 25696
rect 35855 25656 35900 25684
rect 35894 25644 35900 25656
rect 35952 25644 35958 25696
rect 37550 25644 37556 25696
rect 37608 25684 37614 25696
rect 37737 25687 37795 25693
rect 37737 25684 37749 25687
rect 37608 25656 37749 25684
rect 37608 25644 37614 25656
rect 37737 25653 37749 25656
rect 37783 25653 37795 25687
rect 37737 25647 37795 25653
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 13357 25483 13415 25489
rect 13357 25449 13369 25483
rect 13403 25480 13415 25483
rect 13998 25480 14004 25492
rect 13403 25452 14004 25480
rect 13403 25449 13415 25452
rect 13357 25443 13415 25449
rect 13998 25440 14004 25452
rect 14056 25440 14062 25492
rect 14093 25483 14151 25489
rect 14093 25449 14105 25483
rect 14139 25480 14151 25483
rect 14734 25480 14740 25492
rect 14139 25452 14740 25480
rect 14139 25449 14151 25452
rect 14093 25443 14151 25449
rect 14734 25440 14740 25452
rect 14792 25440 14798 25492
rect 15105 25483 15163 25489
rect 15105 25449 15117 25483
rect 15151 25480 15163 25483
rect 15378 25480 15384 25492
rect 15151 25452 15384 25480
rect 15151 25449 15163 25452
rect 15105 25443 15163 25449
rect 15378 25440 15384 25452
rect 15436 25440 15442 25492
rect 15746 25480 15752 25492
rect 15707 25452 15752 25480
rect 15746 25440 15752 25452
rect 15804 25440 15810 25492
rect 17405 25483 17463 25489
rect 17405 25449 17417 25483
rect 17451 25480 17463 25483
rect 18046 25480 18052 25492
rect 17451 25452 18052 25480
rect 17451 25449 17463 25452
rect 17405 25443 17463 25449
rect 18046 25440 18052 25452
rect 18104 25440 18110 25492
rect 20625 25483 20683 25489
rect 20625 25449 20637 25483
rect 20671 25480 20683 25483
rect 21082 25480 21088 25492
rect 20671 25452 21088 25480
rect 20671 25449 20683 25452
rect 20625 25443 20683 25449
rect 21082 25440 21088 25452
rect 21140 25440 21146 25492
rect 22097 25483 22155 25489
rect 22097 25449 22109 25483
rect 22143 25480 22155 25483
rect 24762 25480 24768 25492
rect 22143 25452 24768 25480
rect 22143 25449 22155 25452
rect 22097 25443 22155 25449
rect 24762 25440 24768 25452
rect 24820 25440 24826 25492
rect 24854 25440 24860 25492
rect 24912 25480 24918 25492
rect 30745 25483 30803 25489
rect 24912 25452 27016 25480
rect 24912 25440 24918 25452
rect 20714 25372 20720 25424
rect 20772 25412 20778 25424
rect 21177 25415 21235 25421
rect 21177 25412 21189 25415
rect 20772 25384 21189 25412
rect 20772 25372 20778 25384
rect 21177 25381 21189 25384
rect 21223 25381 21235 25415
rect 21177 25375 21235 25381
rect 22646 25372 22652 25424
rect 22704 25412 22710 25424
rect 22741 25415 22799 25421
rect 22741 25412 22753 25415
rect 22704 25384 22753 25412
rect 22704 25372 22710 25384
rect 22741 25381 22753 25384
rect 22787 25412 22799 25415
rect 23382 25412 23388 25424
rect 22787 25384 23388 25412
rect 22787 25381 22799 25384
rect 22741 25375 22799 25381
rect 23382 25372 23388 25384
rect 23440 25372 23446 25424
rect 23474 25372 23480 25424
rect 23532 25412 23538 25424
rect 25685 25415 25743 25421
rect 25685 25412 25697 25415
rect 23532 25384 25697 25412
rect 23532 25372 23538 25384
rect 25685 25381 25697 25384
rect 25731 25381 25743 25415
rect 26988 25412 27016 25452
rect 30745 25449 30757 25483
rect 30791 25480 30803 25483
rect 31018 25480 31024 25492
rect 30791 25452 31024 25480
rect 30791 25449 30803 25452
rect 30745 25443 30803 25449
rect 31018 25440 31024 25452
rect 31076 25480 31082 25492
rect 31202 25480 31208 25492
rect 31076 25452 31208 25480
rect 31076 25440 31082 25452
rect 31202 25440 31208 25452
rect 31260 25440 31266 25492
rect 34701 25483 34759 25489
rect 34701 25449 34713 25483
rect 34747 25480 34759 25483
rect 34790 25480 34796 25492
rect 34747 25452 34796 25480
rect 34747 25449 34759 25452
rect 34701 25443 34759 25449
rect 34790 25440 34796 25452
rect 34848 25440 34854 25492
rect 35989 25483 36047 25489
rect 35989 25449 36001 25483
rect 36035 25480 36047 25483
rect 36170 25480 36176 25492
rect 36035 25452 36176 25480
rect 36035 25449 36047 25452
rect 35989 25443 36047 25449
rect 36170 25440 36176 25452
rect 36228 25440 36234 25492
rect 28810 25412 28816 25424
rect 26988 25384 28816 25412
rect 25685 25375 25743 25381
rect 15378 25304 15384 25356
rect 15436 25344 15442 25356
rect 16390 25344 16396 25356
rect 15436 25316 16396 25344
rect 15436 25304 15442 25316
rect 16390 25304 16396 25316
rect 16448 25304 16454 25356
rect 21910 25304 21916 25356
rect 21968 25344 21974 25356
rect 22830 25344 22836 25356
rect 21968 25316 22508 25344
rect 22791 25316 22836 25344
rect 21968 25304 21974 25316
rect 13541 25279 13599 25285
rect 13541 25245 13553 25279
rect 13587 25276 13599 25279
rect 14090 25276 14096 25288
rect 13587 25248 14096 25276
rect 13587 25245 13599 25248
rect 13541 25239 13599 25245
rect 14090 25236 14096 25248
rect 14148 25236 14154 25288
rect 14274 25276 14280 25288
rect 14235 25248 14280 25276
rect 14274 25236 14280 25248
rect 14332 25236 14338 25288
rect 15286 25276 15292 25288
rect 15247 25248 15292 25276
rect 15286 25236 15292 25248
rect 15344 25236 15350 25288
rect 15933 25279 15991 25285
rect 15933 25245 15945 25279
rect 15979 25276 15991 25279
rect 16114 25276 16120 25288
rect 15979 25248 16120 25276
rect 15979 25245 15991 25248
rect 15933 25239 15991 25245
rect 16114 25236 16120 25248
rect 16172 25236 16178 25288
rect 16666 25276 16672 25288
rect 16627 25248 16672 25276
rect 16666 25236 16672 25248
rect 16724 25236 16730 25288
rect 17954 25236 17960 25288
rect 18012 25276 18018 25288
rect 18601 25279 18659 25285
rect 18601 25276 18613 25279
rect 18012 25248 18613 25276
rect 18012 25236 18018 25248
rect 18601 25245 18613 25248
rect 18647 25245 18659 25279
rect 18601 25239 18659 25245
rect 19426 25236 19432 25288
rect 19484 25276 19490 25288
rect 19613 25279 19671 25285
rect 19613 25276 19625 25279
rect 19484 25248 19625 25276
rect 19484 25236 19490 25248
rect 19613 25245 19625 25248
rect 19659 25245 19671 25279
rect 19613 25239 19671 25245
rect 19889 25279 19947 25285
rect 19889 25245 19901 25279
rect 19935 25276 19947 25279
rect 20070 25276 20076 25288
rect 19935 25248 20076 25276
rect 19935 25245 19947 25248
rect 19889 25239 19947 25245
rect 20070 25236 20076 25248
rect 20128 25236 20134 25288
rect 20990 25236 20996 25288
rect 21048 25276 21054 25288
rect 22480 25285 22508 25316
rect 22830 25304 22836 25316
rect 22888 25304 22894 25356
rect 23661 25347 23719 25353
rect 23661 25313 23673 25347
rect 23707 25344 23719 25347
rect 23707 25316 23796 25344
rect 23707 25313 23719 25316
rect 23661 25307 23719 25313
rect 23768 25288 23796 25316
rect 23842 25304 23848 25356
rect 23900 25344 23906 25356
rect 23900 25316 23945 25344
rect 23900 25304 23906 25316
rect 25866 25304 25872 25356
rect 25924 25344 25930 25356
rect 27614 25344 27620 25356
rect 25924 25316 27620 25344
rect 25924 25304 25930 25316
rect 27614 25304 27620 25316
rect 27672 25304 27678 25356
rect 21085 25279 21143 25285
rect 21085 25276 21097 25279
rect 21048 25248 21097 25276
rect 21048 25236 21054 25248
rect 21085 25245 21097 25248
rect 21131 25245 21143 25279
rect 21085 25239 21143 25245
rect 22465 25279 22523 25285
rect 22465 25245 22477 25279
rect 22511 25245 22523 25279
rect 22465 25239 22523 25245
rect 22554 25236 22560 25288
rect 22612 25276 22618 25288
rect 23569 25279 23627 25285
rect 22612 25248 22657 25276
rect 22612 25236 22618 25248
rect 23569 25245 23581 25279
rect 23615 25245 23627 25279
rect 23569 25239 23627 25245
rect 21358 25168 21364 25220
rect 21416 25208 21422 25220
rect 23584 25208 23612 25239
rect 23750 25236 23756 25288
rect 23808 25236 23814 25288
rect 24394 25276 24400 25288
rect 24355 25248 24400 25276
rect 24394 25236 24400 25248
rect 24452 25236 24458 25288
rect 24670 25276 24676 25288
rect 24631 25248 24676 25276
rect 24670 25236 24676 25248
rect 24728 25236 24734 25288
rect 25961 25279 26019 25285
rect 25961 25276 25973 25279
rect 24780 25248 25973 25276
rect 21416 25180 23612 25208
rect 21416 25168 21422 25180
rect 24118 25168 24124 25220
rect 24176 25208 24182 25220
rect 24780 25208 24808 25248
rect 25961 25245 25973 25248
rect 26007 25276 26019 25279
rect 26510 25276 26516 25288
rect 26007 25248 26516 25276
rect 26007 25245 26019 25248
rect 25961 25239 26019 25245
rect 26510 25236 26516 25248
rect 26568 25236 26574 25288
rect 26878 25276 26884 25288
rect 26839 25248 26884 25276
rect 26878 25236 26884 25248
rect 26936 25236 26942 25288
rect 27062 25276 27068 25288
rect 27023 25248 27068 25276
rect 27062 25236 27068 25248
rect 27120 25236 27126 25288
rect 24176 25180 24808 25208
rect 25685 25211 25743 25217
rect 24176 25168 24182 25180
rect 25685 25177 25697 25211
rect 25731 25208 25743 25211
rect 26694 25208 26700 25220
rect 25731 25180 26700 25208
rect 25731 25177 25743 25180
rect 25685 25171 25743 25177
rect 26694 25168 26700 25180
rect 26752 25168 26758 25220
rect 28000 25208 28028 25384
rect 28810 25372 28816 25384
rect 28868 25372 28874 25424
rect 29825 25415 29883 25421
rect 29825 25381 29837 25415
rect 29871 25412 29883 25415
rect 30374 25412 30380 25424
rect 29871 25384 30380 25412
rect 29871 25381 29883 25384
rect 29825 25375 29883 25381
rect 30374 25372 30380 25384
rect 30432 25372 30438 25424
rect 31726 25384 33364 25412
rect 28626 25344 28632 25356
rect 28184 25316 28632 25344
rect 28074 25236 28080 25288
rect 28132 25276 28138 25288
rect 28184 25285 28212 25316
rect 28626 25304 28632 25316
rect 28684 25304 28690 25356
rect 30006 25304 30012 25356
rect 30064 25344 30070 25356
rect 30064 25316 31616 25344
rect 30064 25304 30070 25316
rect 28169 25279 28227 25285
rect 28169 25276 28181 25279
rect 28132 25248 28181 25276
rect 28132 25236 28138 25248
rect 28169 25245 28181 25248
rect 28215 25245 28227 25279
rect 28169 25239 28227 25245
rect 28261 25279 28319 25285
rect 28261 25245 28273 25279
rect 28307 25245 28319 25279
rect 28261 25239 28319 25245
rect 28445 25279 28503 25285
rect 28445 25245 28457 25279
rect 28491 25245 28503 25279
rect 28445 25239 28503 25245
rect 28276 25208 28304 25239
rect 28000 25180 28304 25208
rect 28460 25208 28488 25239
rect 28534 25236 28540 25288
rect 28592 25276 28598 25288
rect 28592 25248 28637 25276
rect 28592 25236 28598 25248
rect 29454 25236 29460 25288
rect 29512 25276 29518 25288
rect 30101 25279 30159 25285
rect 30101 25276 30113 25279
rect 29512 25248 30113 25276
rect 29512 25236 29518 25248
rect 30101 25245 30113 25248
rect 30147 25245 30159 25279
rect 30650 25276 30656 25288
rect 30101 25239 30159 25245
rect 30300 25248 30656 25276
rect 29086 25208 29092 25220
rect 28460 25180 29092 25208
rect 29086 25168 29092 25180
rect 29144 25168 29150 25220
rect 29825 25211 29883 25217
rect 29825 25177 29837 25211
rect 29871 25208 29883 25211
rect 30300 25208 30328 25248
rect 30650 25236 30656 25248
rect 30708 25276 30714 25288
rect 31202 25276 31208 25288
rect 30708 25248 31208 25276
rect 30708 25236 30714 25248
rect 31202 25236 31208 25248
rect 31260 25236 31266 25288
rect 31588 25285 31616 25316
rect 31573 25279 31631 25285
rect 31573 25245 31585 25279
rect 31619 25245 31631 25279
rect 31573 25239 31631 25245
rect 29871 25180 30328 25208
rect 30561 25211 30619 25217
rect 29871 25177 29883 25180
rect 29825 25171 29883 25177
rect 30561 25177 30573 25211
rect 30607 25208 30619 25211
rect 31294 25208 31300 25220
rect 30607 25180 31300 25208
rect 30607 25177 30619 25180
rect 30561 25171 30619 25177
rect 31294 25168 31300 25180
rect 31352 25208 31358 25220
rect 31726 25208 31754 25384
rect 33336 25353 33364 25384
rect 33321 25347 33379 25353
rect 33321 25313 33333 25347
rect 33367 25344 33379 25347
rect 34054 25344 34060 25356
rect 33367 25316 34060 25344
rect 33367 25313 33379 25316
rect 33321 25307 33379 25313
rect 34054 25304 34060 25316
rect 34112 25304 34118 25356
rect 34514 25304 34520 25356
rect 34572 25344 34578 25356
rect 35345 25347 35403 25353
rect 35345 25344 35357 25347
rect 34572 25316 35357 25344
rect 34572 25304 34578 25316
rect 35345 25313 35357 25316
rect 35391 25313 35403 25347
rect 37550 25344 37556 25356
rect 37511 25316 37556 25344
rect 35345 25307 35403 25313
rect 37550 25304 37556 25316
rect 37608 25304 37614 25356
rect 32306 25236 32312 25288
rect 32364 25276 32370 25288
rect 32493 25279 32551 25285
rect 32493 25276 32505 25279
rect 32364 25248 32505 25276
rect 32364 25236 32370 25248
rect 32493 25245 32505 25248
rect 32539 25245 32551 25279
rect 32493 25239 32551 25245
rect 32677 25279 32735 25285
rect 32677 25245 32689 25279
rect 32723 25276 32735 25279
rect 32858 25276 32864 25288
rect 32723 25248 32864 25276
rect 32723 25245 32735 25248
rect 32677 25239 32735 25245
rect 31352 25180 31754 25208
rect 32508 25208 32536 25239
rect 32858 25236 32864 25248
rect 32916 25236 32922 25288
rect 33597 25279 33655 25285
rect 33597 25245 33609 25279
rect 33643 25245 33655 25279
rect 34072 25276 34100 25304
rect 34826 25279 34884 25285
rect 34826 25276 34838 25279
rect 34072 25248 34838 25276
rect 33597 25239 33655 25245
rect 34826 25245 34838 25248
rect 34872 25245 34884 25279
rect 35250 25276 35256 25288
rect 35211 25248 35256 25276
rect 34826 25239 34884 25245
rect 33612 25208 33640 25239
rect 35250 25236 35256 25248
rect 35308 25236 35314 25288
rect 37461 25279 37519 25285
rect 37461 25245 37473 25279
rect 37507 25276 37519 25279
rect 37826 25276 37832 25288
rect 37507 25248 37832 25276
rect 37507 25245 37519 25248
rect 37461 25239 37519 25245
rect 37826 25236 37832 25248
rect 37884 25236 37890 25288
rect 35710 25208 35716 25220
rect 32508 25180 35716 25208
rect 31352 25168 31358 25180
rect 18417 25143 18475 25149
rect 18417 25109 18429 25143
rect 18463 25140 18475 25143
rect 18598 25140 18604 25152
rect 18463 25112 18604 25140
rect 18463 25109 18475 25112
rect 18417 25103 18475 25109
rect 18598 25100 18604 25112
rect 18656 25100 18662 25152
rect 22379 25143 22437 25149
rect 22379 25109 22391 25143
rect 22425 25140 22437 25143
rect 23382 25140 23388 25152
rect 22425 25112 23388 25140
rect 22425 25109 22437 25112
rect 22379 25103 22437 25109
rect 23382 25100 23388 25112
rect 23440 25100 23446 25152
rect 23566 25100 23572 25152
rect 23624 25140 23630 25152
rect 23845 25143 23903 25149
rect 23845 25140 23857 25143
rect 23624 25112 23857 25140
rect 23624 25100 23630 25112
rect 23845 25109 23857 25112
rect 23891 25109 23903 25143
rect 25866 25140 25872 25152
rect 25827 25112 25872 25140
rect 23845 25103 23903 25109
rect 25866 25100 25872 25112
rect 25924 25100 25930 25152
rect 26510 25100 26516 25152
rect 26568 25140 26574 25152
rect 26973 25143 27031 25149
rect 26973 25140 26985 25143
rect 26568 25112 26985 25140
rect 26568 25100 26574 25112
rect 26973 25109 26985 25112
rect 27019 25109 27031 25143
rect 26973 25103 27031 25109
rect 27614 25100 27620 25152
rect 27672 25140 27678 25152
rect 27985 25143 28043 25149
rect 27985 25140 27997 25143
rect 27672 25112 27997 25140
rect 27672 25100 27678 25112
rect 27985 25109 27997 25112
rect 28031 25109 28043 25143
rect 27985 25103 28043 25109
rect 30009 25143 30067 25149
rect 30009 25109 30021 25143
rect 30055 25140 30067 25143
rect 30650 25140 30656 25152
rect 30055 25112 30656 25140
rect 30055 25109 30067 25112
rect 30009 25103 30067 25109
rect 30650 25100 30656 25112
rect 30708 25100 30714 25152
rect 30742 25100 30748 25152
rect 30800 25149 30806 25152
rect 30800 25143 30819 25149
rect 30807 25109 30819 25143
rect 30926 25140 30932 25152
rect 30887 25112 30932 25140
rect 30800 25103 30819 25109
rect 30800 25100 30806 25103
rect 30926 25100 30932 25112
rect 30984 25100 30990 25152
rect 31404 25149 31432 25180
rect 35710 25168 35716 25180
rect 35768 25208 35774 25220
rect 35805 25211 35863 25217
rect 35805 25208 35817 25211
rect 35768 25180 35817 25208
rect 35768 25168 35774 25180
rect 35805 25177 35817 25180
rect 35851 25177 35863 25211
rect 35805 25171 35863 25177
rect 31389 25143 31447 25149
rect 31389 25109 31401 25143
rect 31435 25109 31447 25143
rect 31389 25103 31447 25109
rect 32214 25100 32220 25152
rect 32272 25140 32278 25152
rect 32585 25143 32643 25149
rect 32585 25140 32597 25143
rect 32272 25112 32597 25140
rect 32272 25100 32278 25112
rect 32585 25109 32597 25112
rect 32631 25109 32643 25143
rect 32585 25103 32643 25109
rect 33686 25100 33692 25152
rect 33744 25140 33750 25152
rect 34885 25143 34943 25149
rect 34885 25140 34897 25143
rect 33744 25112 34897 25140
rect 33744 25100 33750 25112
rect 34885 25109 34897 25112
rect 34931 25109 34943 25143
rect 34885 25103 34943 25109
rect 35986 25100 35992 25152
rect 36044 25149 36050 25152
rect 36044 25143 36063 25149
rect 36051 25109 36063 25143
rect 36170 25140 36176 25152
rect 36131 25112 36176 25140
rect 36044 25103 36063 25109
rect 36044 25100 36050 25103
rect 36170 25100 36176 25112
rect 36228 25100 36234 25152
rect 37550 25100 37556 25152
rect 37608 25140 37614 25152
rect 37829 25143 37887 25149
rect 37829 25140 37841 25143
rect 37608 25112 37841 25140
rect 37608 25100 37614 25112
rect 37829 25109 37841 25112
rect 37875 25109 37887 25143
rect 37829 25103 37887 25109
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 14274 24896 14280 24948
rect 14332 24936 14338 24948
rect 14553 24939 14611 24945
rect 14553 24936 14565 24939
rect 14332 24908 14565 24936
rect 14332 24896 14338 24908
rect 14553 24905 14565 24908
rect 14599 24905 14611 24939
rect 18966 24936 18972 24948
rect 14553 24899 14611 24905
rect 15028 24908 18972 24936
rect 15028 24880 15056 24908
rect 18966 24896 18972 24908
rect 19024 24896 19030 24948
rect 19058 24896 19064 24948
rect 19116 24936 19122 24948
rect 24302 24936 24308 24948
rect 19116 24908 24308 24936
rect 19116 24896 19122 24908
rect 24302 24896 24308 24908
rect 24360 24896 24366 24948
rect 24394 24896 24400 24948
rect 24452 24936 24458 24948
rect 24581 24939 24639 24945
rect 24581 24936 24593 24939
rect 24452 24908 24593 24936
rect 24452 24896 24458 24908
rect 24581 24905 24593 24908
rect 24627 24905 24639 24939
rect 24581 24899 24639 24905
rect 26234 24896 26240 24948
rect 26292 24936 26298 24948
rect 26421 24939 26479 24945
rect 26421 24936 26433 24939
rect 26292 24908 26433 24936
rect 26292 24896 26298 24908
rect 26421 24905 26433 24908
rect 26467 24905 26479 24939
rect 26421 24899 26479 24905
rect 31570 24896 31576 24948
rect 31628 24936 31634 24948
rect 31938 24936 31944 24948
rect 31628 24908 31944 24936
rect 31628 24896 31634 24908
rect 31938 24896 31944 24908
rect 31996 24936 32002 24948
rect 32861 24939 32919 24945
rect 32861 24936 32873 24939
rect 31996 24908 32873 24936
rect 31996 24896 32002 24908
rect 32861 24905 32873 24908
rect 32907 24905 32919 24939
rect 34054 24936 34060 24948
rect 34015 24908 34060 24936
rect 32861 24899 32919 24905
rect 34054 24896 34060 24908
rect 34112 24896 34118 24948
rect 37277 24939 37335 24945
rect 37277 24905 37289 24939
rect 37323 24936 37335 24939
rect 37458 24936 37464 24948
rect 37323 24908 37464 24936
rect 37323 24905 37335 24908
rect 37277 24899 37335 24905
rect 37458 24896 37464 24908
rect 37516 24896 37522 24948
rect 12986 24828 12992 24880
rect 13044 24868 13050 24880
rect 13357 24871 13415 24877
rect 13357 24868 13369 24871
rect 13044 24840 13369 24868
rect 13044 24828 13050 24840
rect 13357 24837 13369 24840
rect 13403 24837 13415 24871
rect 13557 24871 13615 24877
rect 13557 24868 13569 24871
rect 13357 24831 13415 24837
rect 13556 24837 13569 24868
rect 13603 24837 13615 24871
rect 13556 24831 13615 24837
rect 13556 24800 13584 24831
rect 13814 24828 13820 24880
rect 13872 24868 13878 24880
rect 14185 24871 14243 24877
rect 14185 24868 14197 24871
rect 13872 24840 14197 24868
rect 13872 24828 13878 24840
rect 14185 24837 14197 24840
rect 14231 24837 14243 24871
rect 14385 24871 14443 24877
rect 14385 24868 14397 24871
rect 14185 24831 14243 24837
rect 14384 24837 14397 24868
rect 14431 24837 14443 24871
rect 15010 24868 15016 24880
rect 14923 24840 15016 24868
rect 14384 24831 14443 24837
rect 14274 24800 14280 24812
rect 13556 24772 14280 24800
rect 14274 24760 14280 24772
rect 14332 24800 14338 24812
rect 14384 24800 14412 24831
rect 15010 24828 15016 24840
rect 15068 24828 15074 24880
rect 15213 24871 15271 24877
rect 15213 24868 15225 24871
rect 15212 24837 15225 24868
rect 15259 24837 15271 24871
rect 24670 24868 24676 24880
rect 15212 24831 15271 24837
rect 21468 24840 22140 24868
rect 15212 24800 15240 24831
rect 14332 24772 15516 24800
rect 14332 24760 14338 24772
rect 10042 24692 10048 24744
rect 10100 24732 10106 24744
rect 15010 24732 15016 24744
rect 10100 24704 15016 24732
rect 10100 24692 10106 24704
rect 15010 24692 15016 24704
rect 15068 24692 15074 24744
rect 15194 24692 15200 24744
rect 15252 24732 15258 24744
rect 15488 24732 15516 24772
rect 15930 24760 15936 24812
rect 15988 24800 15994 24812
rect 16117 24803 16175 24809
rect 16117 24800 16129 24803
rect 15988 24772 16129 24800
rect 15988 24760 15994 24772
rect 16117 24769 16129 24772
rect 16163 24769 16175 24803
rect 16117 24763 16175 24769
rect 17129 24803 17187 24809
rect 17129 24769 17141 24803
rect 17175 24800 17187 24803
rect 18046 24800 18052 24812
rect 17175 24772 18052 24800
rect 17175 24769 17187 24772
rect 17129 24763 17187 24769
rect 18046 24760 18052 24772
rect 18104 24760 18110 24812
rect 18598 24800 18604 24812
rect 18559 24772 18604 24800
rect 18598 24760 18604 24772
rect 18656 24760 18662 24812
rect 19794 24760 19800 24812
rect 19852 24800 19858 24812
rect 19981 24803 20039 24809
rect 19981 24800 19993 24803
rect 19852 24772 19993 24800
rect 19852 24760 19858 24772
rect 19981 24769 19993 24772
rect 20027 24769 20039 24803
rect 20438 24800 20444 24812
rect 20399 24772 20444 24800
rect 19981 24763 20039 24769
rect 20438 24760 20444 24772
rect 20496 24760 20502 24812
rect 20530 24760 20536 24812
rect 20588 24800 20594 24812
rect 21085 24803 21143 24809
rect 20588 24772 20633 24800
rect 20588 24760 20594 24772
rect 21085 24769 21097 24803
rect 21131 24800 21143 24803
rect 21174 24800 21180 24812
rect 21131 24772 21180 24800
rect 21131 24769 21143 24772
rect 21085 24763 21143 24769
rect 21174 24760 21180 24772
rect 21232 24760 21238 24812
rect 21266 24760 21272 24812
rect 21324 24800 21330 24812
rect 21324 24772 21369 24800
rect 21324 24760 21330 24772
rect 16758 24732 16764 24744
rect 15252 24704 15424 24732
rect 15488 24704 16764 24732
rect 15252 24692 15258 24704
rect 13725 24667 13783 24673
rect 13725 24633 13737 24667
rect 13771 24664 13783 24667
rect 14642 24664 14648 24676
rect 13771 24636 14648 24664
rect 13771 24633 13783 24636
rect 13725 24627 13783 24633
rect 14642 24624 14648 24636
rect 14700 24624 14706 24676
rect 15396 24673 15424 24704
rect 16758 24692 16764 24704
rect 16816 24692 16822 24744
rect 16853 24735 16911 24741
rect 16853 24701 16865 24735
rect 16899 24701 16911 24735
rect 16853 24695 16911 24701
rect 18325 24735 18383 24741
rect 18325 24701 18337 24735
rect 18371 24701 18383 24735
rect 21468 24732 21496 24840
rect 21726 24760 21732 24812
rect 21784 24800 21790 24812
rect 22112 24809 22140 24840
rect 23400 24840 24676 24868
rect 21821 24803 21879 24809
rect 21821 24800 21833 24803
rect 21784 24772 21833 24800
rect 21784 24760 21790 24772
rect 21821 24769 21833 24772
rect 21867 24769 21879 24803
rect 21821 24763 21879 24769
rect 22097 24803 22155 24809
rect 22097 24769 22109 24803
rect 22143 24769 22155 24803
rect 22097 24763 22155 24769
rect 23014 24760 23020 24812
rect 23072 24800 23078 24812
rect 23400 24809 23428 24840
rect 24670 24828 24676 24840
rect 24728 24828 24734 24880
rect 25222 24828 25228 24880
rect 25280 24868 25286 24880
rect 25409 24871 25467 24877
rect 25409 24868 25421 24871
rect 25280 24840 25421 24868
rect 25280 24828 25286 24840
rect 25409 24837 25421 24840
rect 25455 24868 25467 24871
rect 26050 24868 26056 24880
rect 25455 24840 26056 24868
rect 25455 24837 25467 24840
rect 25409 24831 25467 24837
rect 26050 24828 26056 24840
rect 26108 24828 26114 24880
rect 27522 24868 27528 24880
rect 27172 24840 27528 24868
rect 23385 24803 23443 24809
rect 23385 24800 23397 24803
rect 23072 24772 23397 24800
rect 23072 24760 23078 24772
rect 23385 24769 23397 24772
rect 23431 24769 23443 24803
rect 23385 24763 23443 24769
rect 23842 24760 23848 24812
rect 23900 24800 23906 24812
rect 24397 24803 24455 24809
rect 24397 24800 24409 24803
rect 23900 24772 24409 24800
rect 23900 24760 23906 24772
rect 24397 24769 24409 24772
rect 24443 24769 24455 24803
rect 24397 24763 24455 24769
rect 25498 24760 25504 24812
rect 25556 24800 25562 24812
rect 25593 24803 25651 24809
rect 25593 24800 25605 24803
rect 25556 24772 25605 24800
rect 25556 24760 25562 24772
rect 25593 24769 25605 24772
rect 25639 24769 25651 24803
rect 25593 24763 25651 24769
rect 25685 24803 25743 24809
rect 25685 24769 25697 24803
rect 25731 24800 25743 24803
rect 25958 24800 25964 24812
rect 25731 24772 25964 24800
rect 25731 24769 25743 24772
rect 25685 24763 25743 24769
rect 25958 24760 25964 24772
rect 26016 24760 26022 24812
rect 26145 24803 26203 24809
rect 26145 24769 26157 24803
rect 26191 24800 26203 24803
rect 26234 24800 26240 24812
rect 26191 24772 26240 24800
rect 26191 24769 26203 24772
rect 26145 24763 26203 24769
rect 26234 24760 26240 24772
rect 26292 24760 26298 24812
rect 26786 24760 26792 24812
rect 26844 24800 26850 24812
rect 27172 24809 27200 24840
rect 27522 24828 27528 24840
rect 27580 24868 27586 24880
rect 28258 24868 28264 24880
rect 27580 24840 28264 24868
rect 27580 24828 27586 24840
rect 28258 24828 28264 24840
rect 28316 24828 28322 24880
rect 31018 24868 31024 24880
rect 30576 24840 31024 24868
rect 26973 24803 27031 24809
rect 26973 24800 26985 24803
rect 26844 24772 26985 24800
rect 26844 24760 26850 24772
rect 26973 24769 26985 24772
rect 27019 24769 27031 24803
rect 26973 24763 27031 24769
rect 27157 24803 27215 24809
rect 27157 24769 27169 24803
rect 27203 24769 27215 24803
rect 28074 24800 28080 24812
rect 28035 24772 28080 24800
rect 27157 24763 27215 24769
rect 18325 24695 18383 24701
rect 19812 24704 21496 24732
rect 15381 24667 15439 24673
rect 15381 24633 15393 24667
rect 15427 24633 15439 24667
rect 15381 24627 15439 24633
rect 15933 24667 15991 24673
rect 15933 24633 15945 24667
rect 15979 24664 15991 24667
rect 16666 24664 16672 24676
rect 15979 24636 16672 24664
rect 15979 24633 15991 24636
rect 15933 24627 15991 24633
rect 16666 24624 16672 24636
rect 16724 24624 16730 24676
rect 13541 24599 13599 24605
rect 13541 24565 13553 24599
rect 13587 24596 13599 24599
rect 14369 24599 14427 24605
rect 14369 24596 14381 24599
rect 13587 24568 14381 24596
rect 13587 24565 13599 24568
rect 13541 24559 13599 24565
rect 14369 24565 14381 24568
rect 14415 24596 14427 24599
rect 15194 24596 15200 24608
rect 14415 24568 15200 24596
rect 14415 24565 14427 24568
rect 14369 24559 14427 24565
rect 15194 24556 15200 24568
rect 15252 24556 15258 24608
rect 16868 24596 16896 24695
rect 17865 24667 17923 24673
rect 17865 24633 17877 24667
rect 17911 24664 17923 24667
rect 18138 24664 18144 24676
rect 17911 24636 18144 24664
rect 17911 24633 17923 24636
rect 17865 24627 17923 24633
rect 18138 24624 18144 24636
rect 18196 24624 18202 24676
rect 17770 24596 17776 24608
rect 16868 24568 17776 24596
rect 17770 24556 17776 24568
rect 17828 24596 17834 24608
rect 18340 24596 18368 24695
rect 19426 24664 19432 24676
rect 19260 24636 19432 24664
rect 19260 24596 19288 24636
rect 19426 24624 19432 24636
rect 19484 24624 19490 24676
rect 19812 24673 19840 24704
rect 22554 24692 22560 24744
rect 22612 24732 22618 24744
rect 23661 24735 23719 24741
rect 23661 24732 23673 24735
rect 22612 24704 23673 24732
rect 22612 24692 22618 24704
rect 23661 24701 23673 24704
rect 23707 24701 23719 24735
rect 23661 24695 23719 24701
rect 24213 24735 24271 24741
rect 24213 24701 24225 24735
rect 24259 24732 24271 24735
rect 24854 24732 24860 24744
rect 24259 24704 24860 24732
rect 24259 24701 24271 24704
rect 24213 24695 24271 24701
rect 24854 24692 24860 24704
rect 24912 24732 24918 24744
rect 25866 24732 25872 24744
rect 24912 24704 25872 24732
rect 24912 24692 24918 24704
rect 25866 24692 25872 24704
rect 25924 24692 25930 24744
rect 26418 24732 26424 24744
rect 26379 24704 26424 24732
rect 26418 24692 26424 24704
rect 26476 24692 26482 24744
rect 26988 24732 27016 24763
rect 28074 24760 28080 24772
rect 28132 24760 28138 24812
rect 28902 24800 28908 24812
rect 28815 24772 28908 24800
rect 28902 24760 28908 24772
rect 28960 24800 28966 24812
rect 30576 24809 30604 24840
rect 31018 24828 31024 24840
rect 31076 24828 31082 24880
rect 31294 24828 31300 24880
rect 31352 24868 31358 24880
rect 33134 24868 33140 24880
rect 31352 24840 32260 24868
rect 31352 24828 31358 24840
rect 30561 24803 30619 24809
rect 28960 24772 30512 24800
rect 28960 24760 28966 24772
rect 27246 24732 27252 24744
rect 26988 24704 27252 24732
rect 27246 24692 27252 24704
rect 27304 24692 27310 24744
rect 30374 24732 30380 24744
rect 30335 24704 30380 24732
rect 30374 24692 30380 24704
rect 30432 24692 30438 24744
rect 30484 24732 30512 24772
rect 30561 24769 30573 24803
rect 30607 24769 30619 24803
rect 30561 24763 30619 24769
rect 30650 24760 30656 24812
rect 30708 24800 30714 24812
rect 30708 24772 31708 24800
rect 30708 24760 30714 24772
rect 30745 24735 30803 24741
rect 30745 24732 30757 24735
rect 30484 24704 30757 24732
rect 30745 24701 30757 24704
rect 30791 24701 30803 24735
rect 31202 24732 31208 24744
rect 31163 24704 31208 24732
rect 30745 24695 30803 24701
rect 31202 24692 31208 24704
rect 31260 24692 31266 24744
rect 31680 24732 31708 24772
rect 32030 24760 32036 24812
rect 32088 24800 32094 24812
rect 32125 24803 32183 24809
rect 32125 24800 32137 24803
rect 32088 24772 32137 24800
rect 32088 24760 32094 24772
rect 32125 24769 32137 24772
rect 32171 24769 32183 24803
rect 32125 24763 32183 24769
rect 32232 24732 32260 24840
rect 32508 24840 33140 24868
rect 32309 24803 32367 24809
rect 32309 24769 32321 24803
rect 32355 24800 32367 24803
rect 32508 24800 32536 24840
rect 33134 24828 33140 24840
rect 33192 24828 33198 24880
rect 34977 24871 35035 24877
rect 34977 24868 34989 24871
rect 33888 24840 34989 24868
rect 33888 24812 33916 24840
rect 34977 24837 34989 24840
rect 35023 24868 35035 24871
rect 35250 24868 35256 24880
rect 35023 24840 35256 24868
rect 35023 24837 35035 24840
rect 34977 24831 35035 24837
rect 35250 24828 35256 24840
rect 35308 24828 35314 24880
rect 35894 24868 35900 24880
rect 35855 24840 35900 24868
rect 35894 24828 35900 24840
rect 35952 24828 35958 24880
rect 32766 24800 32772 24812
rect 32355 24772 32536 24800
rect 32727 24772 32772 24800
rect 32355 24769 32367 24772
rect 32309 24763 32367 24769
rect 32766 24760 32772 24772
rect 32824 24760 32830 24812
rect 32953 24803 33011 24809
rect 32953 24769 32965 24803
rect 32999 24769 33011 24803
rect 32953 24763 33011 24769
rect 33689 24803 33747 24809
rect 33689 24769 33701 24803
rect 33735 24800 33747 24803
rect 33870 24800 33876 24812
rect 33735 24772 33876 24800
rect 33735 24769 33747 24772
rect 33689 24763 33747 24769
rect 32968 24732 32996 24763
rect 33870 24760 33876 24772
rect 33928 24760 33934 24812
rect 34174 24803 34232 24809
rect 34174 24769 34186 24803
rect 34220 24800 34232 24803
rect 34330 24800 34336 24812
rect 34220 24772 34336 24800
rect 34220 24769 34232 24772
rect 34174 24763 34232 24769
rect 34330 24760 34336 24772
rect 34388 24760 34394 24812
rect 34811 24803 34869 24809
rect 34811 24769 34823 24803
rect 34857 24769 34869 24803
rect 34811 24763 34869 24769
rect 35161 24803 35219 24809
rect 35161 24769 35173 24803
rect 35207 24800 35219 24803
rect 35986 24800 35992 24812
rect 35207 24772 35992 24800
rect 35207 24769 35219 24772
rect 35161 24763 35219 24769
rect 31680 24704 32168 24732
rect 32232 24704 32996 24732
rect 19797 24667 19855 24673
rect 19797 24633 19809 24667
rect 19843 24633 19855 24667
rect 19797 24627 19855 24633
rect 21266 24624 21272 24676
rect 21324 24664 21330 24676
rect 23474 24664 23480 24676
rect 21324 24636 21956 24664
rect 23435 24636 23480 24664
rect 21324 24624 21330 24636
rect 17828 24568 19288 24596
rect 19337 24599 19395 24605
rect 17828 24556 17834 24568
rect 19337 24565 19349 24599
rect 19383 24596 19395 24599
rect 20714 24596 20720 24608
rect 19383 24568 20720 24596
rect 19383 24565 19395 24568
rect 19337 24559 19395 24565
rect 20714 24556 20720 24568
rect 20772 24556 20778 24608
rect 21177 24599 21235 24605
rect 21177 24565 21189 24599
rect 21223 24596 21235 24599
rect 21818 24596 21824 24608
rect 21223 24568 21824 24596
rect 21223 24565 21235 24568
rect 21177 24559 21235 24565
rect 21818 24556 21824 24568
rect 21876 24556 21882 24608
rect 21928 24596 21956 24636
rect 23474 24624 23480 24636
rect 23532 24624 23538 24676
rect 29270 24664 29276 24676
rect 29231 24636 29276 24664
rect 29270 24624 29276 24636
rect 29328 24624 29334 24676
rect 31113 24667 31171 24673
rect 31113 24633 31125 24667
rect 31159 24664 31171 24667
rect 32030 24664 32036 24676
rect 31159 24636 32036 24664
rect 31159 24633 31171 24636
rect 31113 24627 31171 24633
rect 32030 24624 32036 24636
rect 32088 24624 32094 24676
rect 32140 24664 32168 24704
rect 33778 24692 33784 24744
rect 33836 24732 33842 24744
rect 33965 24735 34023 24741
rect 33965 24732 33977 24735
rect 33836 24704 33977 24732
rect 33836 24692 33842 24704
rect 33965 24701 33977 24704
rect 34011 24701 34023 24735
rect 33965 24695 34023 24701
rect 34841 24676 34869 24763
rect 35986 24760 35992 24772
rect 36044 24760 36050 24812
rect 36081 24803 36139 24809
rect 36081 24769 36093 24803
rect 36127 24769 36139 24803
rect 36081 24763 36139 24769
rect 36096 24732 36124 24763
rect 36722 24760 36728 24812
rect 36780 24800 36786 24812
rect 37461 24803 37519 24809
rect 37461 24800 37473 24803
rect 36780 24772 37473 24800
rect 36780 24760 36786 24772
rect 37461 24769 37473 24772
rect 37507 24769 37519 24803
rect 37461 24763 37519 24769
rect 37645 24803 37703 24809
rect 37645 24769 37657 24803
rect 37691 24769 37703 24803
rect 37645 24763 37703 24769
rect 36170 24732 36176 24744
rect 36083 24704 36176 24732
rect 36170 24692 36176 24704
rect 36228 24732 36234 24744
rect 37182 24732 37188 24744
rect 36228 24704 37188 24732
rect 36228 24692 36234 24704
rect 37182 24692 37188 24704
rect 37240 24732 37246 24744
rect 37660 24732 37688 24763
rect 37734 24760 37740 24812
rect 37792 24800 37798 24812
rect 37792 24772 37837 24800
rect 37792 24760 37798 24772
rect 37240 24704 37688 24732
rect 37240 24692 37246 24704
rect 32217 24667 32275 24673
rect 32217 24664 32229 24667
rect 32140 24636 32229 24664
rect 32217 24633 32229 24636
rect 32263 24664 32275 24667
rect 32766 24664 32772 24676
rect 32263 24636 32772 24664
rect 32263 24633 32275 24636
rect 32217 24627 32275 24633
rect 32766 24624 32772 24636
rect 32824 24624 32830 24676
rect 34333 24667 34391 24673
rect 34333 24633 34345 24667
rect 34379 24664 34391 24667
rect 34790 24664 34796 24676
rect 34379 24636 34796 24664
rect 34379 24633 34391 24636
rect 34333 24627 34391 24633
rect 34790 24624 34796 24636
rect 34848 24636 34869 24676
rect 34848 24624 34854 24636
rect 22738 24596 22744 24608
rect 21928 24568 22744 24596
rect 22738 24556 22744 24568
rect 22796 24556 22802 24608
rect 22833 24599 22891 24605
rect 22833 24565 22845 24599
rect 22879 24596 22891 24599
rect 23106 24596 23112 24608
rect 22879 24568 23112 24596
rect 22879 24565 22891 24568
rect 22833 24559 22891 24565
rect 23106 24556 23112 24568
rect 23164 24556 23170 24608
rect 23569 24599 23627 24605
rect 23569 24565 23581 24599
rect 23615 24596 23627 24599
rect 23658 24596 23664 24608
rect 23615 24568 23664 24596
rect 23615 24565 23627 24568
rect 23569 24559 23627 24565
rect 23658 24556 23664 24568
rect 23716 24556 23722 24608
rect 23750 24556 23756 24608
rect 23808 24596 23814 24608
rect 25409 24599 25467 24605
rect 25409 24596 25421 24599
rect 23808 24568 25421 24596
rect 23808 24556 23814 24568
rect 25409 24565 25421 24568
rect 25455 24565 25467 24599
rect 26234 24596 26240 24608
rect 26195 24568 26240 24596
rect 25409 24559 25467 24565
rect 26234 24556 26240 24568
rect 26292 24556 26298 24608
rect 26786 24556 26792 24608
rect 26844 24596 26850 24608
rect 27062 24596 27068 24608
rect 26844 24568 27068 24596
rect 26844 24556 26850 24568
rect 27062 24556 27068 24568
rect 27120 24596 27126 24608
rect 27341 24599 27399 24605
rect 27341 24596 27353 24599
rect 27120 24568 27353 24596
rect 27120 24556 27126 24568
rect 27341 24565 27353 24568
rect 27387 24565 27399 24599
rect 27341 24559 27399 24565
rect 31570 24556 31576 24608
rect 31628 24596 31634 24608
rect 31846 24596 31852 24608
rect 31628 24568 31852 24596
rect 31628 24556 31634 24568
rect 31846 24556 31852 24568
rect 31904 24556 31910 24608
rect 32398 24556 32404 24608
rect 32456 24596 32462 24608
rect 35434 24596 35440 24608
rect 32456 24568 35440 24596
rect 32456 24556 32462 24568
rect 35434 24556 35440 24568
rect 35492 24556 35498 24608
rect 36262 24596 36268 24608
rect 36223 24568 36268 24596
rect 36262 24556 36268 24568
rect 36320 24556 36326 24608
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 14277 24395 14335 24401
rect 14277 24361 14289 24395
rect 14323 24392 14335 24395
rect 15105 24395 15163 24401
rect 14323 24364 14872 24392
rect 14323 24361 14335 24364
rect 14277 24355 14335 24361
rect 13906 24284 13912 24336
rect 13964 24324 13970 24336
rect 14461 24327 14519 24333
rect 14461 24324 14473 24327
rect 13964 24296 14473 24324
rect 13964 24284 13970 24296
rect 14461 24293 14473 24296
rect 14507 24293 14519 24327
rect 14844 24324 14872 24364
rect 15105 24361 15117 24395
rect 15151 24392 15163 24395
rect 15933 24395 15991 24401
rect 15933 24392 15945 24395
rect 15151 24364 15945 24392
rect 15151 24361 15163 24364
rect 15105 24355 15163 24361
rect 15933 24361 15945 24364
rect 15979 24361 15991 24395
rect 16114 24392 16120 24404
rect 16075 24364 16120 24392
rect 15933 24355 15991 24361
rect 15194 24324 15200 24336
rect 14844 24296 15200 24324
rect 14461 24287 14519 24293
rect 15194 24284 15200 24296
rect 15252 24284 15258 24336
rect 15286 24284 15292 24336
rect 15344 24324 15350 24336
rect 15948 24324 15976 24355
rect 16114 24352 16120 24364
rect 16172 24352 16178 24404
rect 16482 24352 16488 24404
rect 16540 24392 16546 24404
rect 16761 24395 16819 24401
rect 16761 24392 16773 24395
rect 16540 24364 16773 24392
rect 16540 24352 16546 24364
rect 16761 24361 16773 24364
rect 16807 24361 16819 24395
rect 16761 24355 16819 24361
rect 19426 24352 19432 24404
rect 19484 24352 19490 24404
rect 19794 24392 19800 24404
rect 19755 24364 19800 24392
rect 19794 24352 19800 24364
rect 19852 24352 19858 24404
rect 20438 24352 20444 24404
rect 20496 24392 20502 24404
rect 20496 24364 22140 24392
rect 20496 24352 20502 24364
rect 16500 24324 16528 24352
rect 15344 24296 15389 24324
rect 15948 24296 16528 24324
rect 16945 24327 17003 24333
rect 15344 24284 15350 24296
rect 16945 24293 16957 24327
rect 16991 24293 17003 24327
rect 19444 24324 19472 24352
rect 22005 24327 22063 24333
rect 19444 24296 21036 24324
rect 16945 24287 17003 24293
rect 10226 24216 10232 24268
rect 10284 24256 10290 24268
rect 11517 24259 11575 24265
rect 11517 24256 11529 24259
rect 10284 24228 11529 24256
rect 10284 24216 10290 24228
rect 11517 24225 11529 24228
rect 11563 24225 11575 24259
rect 11517 24219 11575 24225
rect 11977 24259 12035 24265
rect 11977 24225 11989 24259
rect 12023 24256 12035 24259
rect 12529 24259 12587 24265
rect 12529 24256 12541 24259
rect 12023 24228 12541 24256
rect 12023 24225 12035 24228
rect 11977 24219 12035 24225
rect 12529 24225 12541 24228
rect 12575 24225 12587 24259
rect 12529 24219 12587 24225
rect 14090 24216 14096 24268
rect 14148 24256 14154 24268
rect 16960 24256 16988 24287
rect 14148 24228 16988 24256
rect 19429 24259 19487 24265
rect 14148 24216 14154 24228
rect 19429 24225 19441 24259
rect 19475 24256 19487 24259
rect 20162 24256 20168 24268
rect 19475 24228 20168 24256
rect 19475 24225 19487 24228
rect 19429 24219 19487 24225
rect 20162 24216 20168 24228
rect 20220 24216 20226 24268
rect 20438 24216 20444 24268
rect 20496 24216 20502 24268
rect 11606 24188 11612 24200
rect 11567 24160 11612 24188
rect 11606 24148 11612 24160
rect 11664 24148 11670 24200
rect 11882 24148 11888 24200
rect 11940 24188 11946 24200
rect 12621 24191 12679 24197
rect 12621 24188 12633 24191
rect 11940 24160 12633 24188
rect 11940 24148 11946 24160
rect 12621 24157 12633 24160
rect 12667 24157 12679 24191
rect 17494 24188 17500 24200
rect 12621 24151 12679 24157
rect 14108 24160 17500 24188
rect 10318 24080 10324 24132
rect 10376 24120 10382 24132
rect 14108 24129 14136 24160
rect 17494 24148 17500 24160
rect 17552 24148 17558 24200
rect 17681 24191 17739 24197
rect 17681 24157 17693 24191
rect 17727 24188 17739 24191
rect 18506 24188 18512 24200
rect 17727 24160 18368 24188
rect 18467 24160 18512 24188
rect 17727 24157 17739 24160
rect 17681 24151 17739 24157
rect 14093 24123 14151 24129
rect 14093 24120 14105 24123
rect 10376 24092 14105 24120
rect 10376 24080 10382 24092
rect 14093 24089 14105 24092
rect 14139 24089 14151 24123
rect 14093 24083 14151 24089
rect 14274 24080 14280 24132
rect 14332 24129 14338 24132
rect 14332 24123 14356 24129
rect 14344 24089 14356 24123
rect 14332 24083 14356 24089
rect 14921 24123 14979 24129
rect 14921 24089 14933 24123
rect 14967 24120 14979 24123
rect 15010 24120 15016 24132
rect 14967 24092 15016 24120
rect 14967 24089 14979 24092
rect 14921 24083 14979 24089
rect 14332 24080 14338 24083
rect 15010 24080 15016 24092
rect 15068 24080 15074 24132
rect 15654 24080 15660 24132
rect 15712 24120 15718 24132
rect 15749 24123 15807 24129
rect 15749 24120 15761 24123
rect 15712 24092 15761 24120
rect 15712 24080 15718 24092
rect 15749 24089 15761 24092
rect 15795 24089 15807 24123
rect 15749 24083 15807 24089
rect 15838 24080 15844 24132
rect 15896 24120 15902 24132
rect 16577 24123 16635 24129
rect 16577 24120 16589 24123
rect 15896 24092 16589 24120
rect 15896 24080 15902 24092
rect 16577 24089 16589 24092
rect 16623 24089 16635 24123
rect 16577 24083 16635 24089
rect 16758 24080 16764 24132
rect 16816 24129 16822 24132
rect 16816 24123 16835 24129
rect 16823 24089 16835 24123
rect 16816 24083 16835 24089
rect 16816 24080 16822 24083
rect 12989 24055 13047 24061
rect 12989 24021 13001 24055
rect 13035 24052 13047 24055
rect 13446 24052 13452 24064
rect 13035 24024 13452 24052
rect 13035 24021 13047 24024
rect 12989 24015 13047 24021
rect 13446 24012 13452 24024
rect 13504 24012 13510 24064
rect 14458 24012 14464 24064
rect 14516 24052 14522 24064
rect 15102 24052 15108 24064
rect 15160 24061 15166 24064
rect 15160 24055 15179 24061
rect 14516 24024 15108 24052
rect 14516 24012 14522 24024
rect 15102 24012 15108 24024
rect 15167 24052 15179 24055
rect 15949 24055 16007 24061
rect 15949 24052 15961 24055
rect 15167 24024 15961 24052
rect 15167 24021 15179 24024
rect 15160 24015 15179 24021
rect 15949 24021 15961 24024
rect 15995 24021 16007 24055
rect 15949 24015 16007 24021
rect 17865 24055 17923 24061
rect 17865 24021 17877 24055
rect 17911 24052 17923 24055
rect 18230 24052 18236 24064
rect 17911 24024 18236 24052
rect 17911 24021 17923 24024
rect 17865 24015 17923 24021
rect 15160 24012 15166 24015
rect 18230 24012 18236 24024
rect 18288 24012 18294 24064
rect 18340 24061 18368 24160
rect 18506 24148 18512 24160
rect 18564 24148 18570 24200
rect 19613 24191 19671 24197
rect 19613 24157 19625 24191
rect 19659 24157 19671 24191
rect 19613 24151 19671 24157
rect 20349 24191 20407 24197
rect 20349 24157 20361 24191
rect 20395 24188 20407 24191
rect 20456 24188 20484 24216
rect 21008 24200 21036 24296
rect 22005 24293 22017 24327
rect 22051 24293 22063 24327
rect 22112 24324 22140 24364
rect 22186 24352 22192 24404
rect 22244 24392 22250 24404
rect 26234 24392 26240 24404
rect 22244 24364 26240 24392
rect 22244 24352 22250 24364
rect 26234 24352 26240 24364
rect 26292 24352 26298 24404
rect 26878 24352 26884 24404
rect 26936 24392 26942 24404
rect 27525 24395 27583 24401
rect 27525 24392 27537 24395
rect 26936 24364 27537 24392
rect 26936 24352 26942 24364
rect 27525 24361 27537 24364
rect 27571 24361 27583 24395
rect 30469 24395 30527 24401
rect 27525 24355 27583 24361
rect 27724 24364 30420 24392
rect 27430 24324 27436 24336
rect 22112 24296 27436 24324
rect 22005 24287 22063 24293
rect 22020 24256 22048 24287
rect 27430 24284 27436 24296
rect 27488 24284 27494 24336
rect 22370 24256 22376 24268
rect 22020 24228 22376 24256
rect 22370 24216 22376 24228
rect 22428 24216 22434 24268
rect 23293 24259 23351 24265
rect 23293 24225 23305 24259
rect 23339 24256 23351 24259
rect 23474 24256 23480 24268
rect 23339 24228 23480 24256
rect 23339 24225 23351 24228
rect 23293 24219 23351 24225
rect 23474 24216 23480 24228
rect 23532 24216 23538 24268
rect 24118 24216 24124 24268
rect 24176 24256 24182 24268
rect 24581 24259 24639 24265
rect 24176 24228 24532 24256
rect 24176 24216 24182 24228
rect 20395 24160 20484 24188
rect 20533 24191 20591 24197
rect 20395 24157 20407 24160
rect 20349 24151 20407 24157
rect 20533 24157 20545 24191
rect 20579 24157 20591 24191
rect 20990 24188 20996 24200
rect 20903 24160 20996 24188
rect 20533 24151 20591 24157
rect 19628 24120 19656 24151
rect 20438 24120 20444 24132
rect 19444 24092 19656 24120
rect 20399 24092 20444 24120
rect 19444 24064 19472 24092
rect 20438 24080 20444 24092
rect 20496 24080 20502 24132
rect 18325 24055 18383 24061
rect 18325 24021 18337 24055
rect 18371 24052 18383 24055
rect 19426 24052 19432 24064
rect 18371 24024 19432 24052
rect 18371 24021 18383 24024
rect 18325 24015 18383 24021
rect 19426 24012 19432 24024
rect 19484 24012 19490 24064
rect 20548 24052 20576 24151
rect 20990 24148 20996 24160
rect 21048 24148 21054 24200
rect 21269 24191 21327 24197
rect 21269 24157 21281 24191
rect 21315 24188 21327 24191
rect 21818 24188 21824 24200
rect 21315 24160 21824 24188
rect 21315 24157 21327 24160
rect 21269 24151 21327 24157
rect 21818 24148 21824 24160
rect 21876 24148 21882 24200
rect 24504 24197 24532 24228
rect 24581 24225 24593 24259
rect 24627 24256 24639 24259
rect 25222 24256 25228 24268
rect 24627 24228 25228 24256
rect 24627 24225 24639 24228
rect 24581 24219 24639 24225
rect 23201 24191 23259 24197
rect 23201 24157 23213 24191
rect 23247 24157 23259 24191
rect 23201 24151 23259 24157
rect 24489 24191 24547 24197
rect 24489 24157 24501 24191
rect 24535 24157 24547 24191
rect 24670 24188 24676 24200
rect 24631 24160 24676 24188
rect 24489 24151 24547 24157
rect 20714 24080 20720 24132
rect 20772 24120 20778 24132
rect 22094 24120 22100 24132
rect 20772 24092 22100 24120
rect 20772 24080 20778 24092
rect 22094 24080 22100 24092
rect 22152 24080 22158 24132
rect 23014 24052 23020 24064
rect 20548 24024 23020 24052
rect 23014 24012 23020 24024
rect 23072 24052 23078 24064
rect 23216 24052 23244 24151
rect 24670 24148 24676 24160
rect 24728 24148 24734 24200
rect 25148 24197 25176 24228
rect 25222 24216 25228 24228
rect 25280 24216 25286 24268
rect 27246 24216 27252 24268
rect 27304 24256 27310 24268
rect 27724 24256 27752 24364
rect 27982 24284 27988 24336
rect 28040 24324 28046 24336
rect 30392 24324 30420 24364
rect 30469 24361 30481 24395
rect 30515 24392 30527 24395
rect 30834 24392 30840 24404
rect 30515 24364 30840 24392
rect 30515 24361 30527 24364
rect 30469 24355 30527 24361
rect 30834 24352 30840 24364
rect 30892 24352 30898 24404
rect 36722 24392 36728 24404
rect 36683 24364 36728 24392
rect 36722 24352 36728 24364
rect 36780 24352 36786 24404
rect 32674 24324 32680 24336
rect 28040 24296 30052 24324
rect 30392 24296 32680 24324
rect 28040 24284 28046 24296
rect 27304 24228 27752 24256
rect 27304 24216 27310 24228
rect 25133 24191 25191 24197
rect 25133 24157 25145 24191
rect 25179 24157 25191 24191
rect 25133 24151 25191 24157
rect 25317 24191 25375 24197
rect 25317 24157 25329 24191
rect 25363 24157 25375 24191
rect 25317 24151 25375 24157
rect 25332 24120 25360 24151
rect 25498 24148 25504 24200
rect 25556 24188 25562 24200
rect 25777 24191 25835 24197
rect 25777 24188 25789 24191
rect 25556 24160 25789 24188
rect 25556 24148 25562 24160
rect 25777 24157 25789 24160
rect 25823 24157 25835 24191
rect 26786 24188 26792 24200
rect 26747 24160 26792 24188
rect 25777 24151 25835 24157
rect 26786 24148 26792 24160
rect 26844 24148 26850 24200
rect 27065 24191 27123 24197
rect 27065 24157 27077 24191
rect 27111 24188 27123 24191
rect 27154 24188 27160 24200
rect 27111 24160 27160 24188
rect 27111 24157 27123 24160
rect 27065 24151 27123 24157
rect 27154 24148 27160 24160
rect 27212 24148 27218 24200
rect 27522 24188 27528 24200
rect 27483 24160 27528 24188
rect 27522 24148 27528 24160
rect 27580 24148 27586 24200
rect 27724 24197 27752 24228
rect 28736 24228 29684 24256
rect 28736 24197 28764 24228
rect 29656 24200 29684 24228
rect 27709 24191 27767 24197
rect 27709 24157 27721 24191
rect 27755 24157 27767 24191
rect 27709 24151 27767 24157
rect 28721 24191 28779 24197
rect 28721 24157 28733 24191
rect 28767 24157 28779 24191
rect 28721 24151 28779 24157
rect 28810 24148 28816 24200
rect 28868 24188 28874 24200
rect 28905 24191 28963 24197
rect 28905 24188 28917 24191
rect 28868 24160 28917 24188
rect 28868 24148 28874 24160
rect 28905 24157 28917 24160
rect 28951 24188 28963 24191
rect 29549 24191 29607 24197
rect 29549 24188 29561 24191
rect 28951 24160 29561 24188
rect 28951 24157 28963 24160
rect 28905 24151 28963 24157
rect 29549 24157 29561 24160
rect 29595 24157 29607 24191
rect 29549 24151 29607 24157
rect 29638 24148 29644 24200
rect 29696 24188 29702 24200
rect 29733 24191 29791 24197
rect 29733 24188 29745 24191
rect 29696 24160 29745 24188
rect 29696 24148 29702 24160
rect 29733 24157 29745 24160
rect 29779 24157 29791 24191
rect 29733 24151 29791 24157
rect 25869 24123 25927 24129
rect 25869 24120 25881 24123
rect 25332 24092 25881 24120
rect 25869 24089 25881 24092
rect 25915 24089 25927 24123
rect 25869 24083 25927 24089
rect 26418 24080 26424 24132
rect 26476 24120 26482 24132
rect 26973 24123 27031 24129
rect 26973 24120 26985 24123
rect 26476 24092 26985 24120
rect 26476 24080 26482 24092
rect 26973 24089 26985 24092
rect 27019 24089 27031 24123
rect 26973 24083 27031 24089
rect 28534 24080 28540 24132
rect 28592 24120 28598 24132
rect 29917 24123 29975 24129
rect 29917 24120 29929 24123
rect 28592 24092 29929 24120
rect 28592 24080 28598 24092
rect 29917 24089 29929 24092
rect 29963 24089 29975 24123
rect 30024 24120 30052 24296
rect 32674 24284 32680 24296
rect 32732 24284 32738 24336
rect 32490 24256 32496 24268
rect 32451 24228 32496 24256
rect 32490 24216 32496 24228
rect 32548 24216 32554 24268
rect 32953 24259 33011 24265
rect 32953 24225 32965 24259
rect 32999 24256 33011 24259
rect 33134 24256 33140 24268
rect 32999 24228 33140 24256
rect 32999 24225 33011 24228
rect 32953 24219 33011 24225
rect 33134 24216 33140 24228
rect 33192 24216 33198 24268
rect 36357 24259 36415 24265
rect 36357 24225 36369 24259
rect 36403 24256 36415 24259
rect 37274 24256 37280 24268
rect 36403 24228 36952 24256
rect 37235 24228 37280 24256
rect 36403 24225 36415 24228
rect 36357 24219 36415 24225
rect 30377 24191 30435 24197
rect 30377 24157 30389 24191
rect 30423 24188 30435 24191
rect 30650 24188 30656 24200
rect 30423 24160 30656 24188
rect 30423 24157 30435 24160
rect 30377 24151 30435 24157
rect 30650 24148 30656 24160
rect 30708 24148 30714 24200
rect 31018 24148 31024 24200
rect 31076 24188 31082 24200
rect 31205 24191 31263 24197
rect 31205 24188 31217 24191
rect 31076 24160 31217 24188
rect 31076 24148 31082 24160
rect 31205 24157 31217 24160
rect 31251 24157 31263 24191
rect 31205 24151 31263 24157
rect 31389 24191 31447 24197
rect 31389 24157 31401 24191
rect 31435 24188 31447 24191
rect 32214 24188 32220 24200
rect 31435 24160 32076 24188
rect 32175 24160 32220 24188
rect 31435 24157 31447 24160
rect 31389 24151 31447 24157
rect 32048 24120 32076 24160
rect 32214 24148 32220 24160
rect 32272 24148 32278 24200
rect 32306 24148 32312 24200
rect 32364 24188 32370 24200
rect 33226 24188 33232 24200
rect 32364 24160 32409 24188
rect 33139 24160 33232 24188
rect 32364 24148 32370 24160
rect 33226 24148 33232 24160
rect 33284 24148 33290 24200
rect 34698 24188 34704 24200
rect 34659 24160 34704 24188
rect 34698 24148 34704 24160
rect 34756 24148 34762 24200
rect 34790 24148 34796 24200
rect 34848 24188 34854 24200
rect 34885 24191 34943 24197
rect 34885 24188 34897 24191
rect 34848 24160 34897 24188
rect 34848 24148 34854 24160
rect 34885 24157 34897 24160
rect 34931 24157 34943 24191
rect 35342 24188 35348 24200
rect 35303 24160 35348 24188
rect 34885 24151 34943 24157
rect 35342 24148 35348 24160
rect 35400 24148 35406 24200
rect 35529 24191 35587 24197
rect 35529 24157 35541 24191
rect 35575 24157 35587 24191
rect 35529 24151 35587 24157
rect 36541 24191 36599 24197
rect 36541 24157 36553 24191
rect 36587 24157 36599 24191
rect 36924 24188 36952 24228
rect 37274 24216 37280 24228
rect 37332 24216 37338 24268
rect 37090 24188 37096 24200
rect 36924 24160 37096 24188
rect 36541 24151 36599 24157
rect 33244 24120 33272 24148
rect 35544 24120 35572 24151
rect 30024 24092 31754 24120
rect 32048 24092 33272 24120
rect 34808 24092 35572 24120
rect 36556 24120 36584 24151
rect 37090 24148 37096 24160
rect 37148 24188 37154 24200
rect 37369 24191 37427 24197
rect 37369 24188 37381 24191
rect 37148 24160 37381 24188
rect 37148 24148 37154 24160
rect 37369 24157 37381 24160
rect 37415 24157 37427 24191
rect 37369 24151 37427 24157
rect 37274 24120 37280 24132
rect 36556 24092 37280 24120
rect 29917 24083 29975 24089
rect 23474 24052 23480 24064
rect 23072 24024 23480 24052
rect 23072 24012 23078 24024
rect 23474 24012 23480 24024
rect 23532 24012 23538 24064
rect 23569 24055 23627 24061
rect 23569 24021 23581 24055
rect 23615 24052 23627 24055
rect 24210 24052 24216 24064
rect 23615 24024 24216 24052
rect 23615 24021 23627 24024
rect 23569 24015 23627 24021
rect 24210 24012 24216 24024
rect 24268 24012 24274 24064
rect 24302 24012 24308 24064
rect 24360 24052 24366 24064
rect 25225 24055 25283 24061
rect 25225 24052 25237 24055
rect 24360 24024 25237 24052
rect 24360 24012 24366 24024
rect 25225 24021 25237 24024
rect 25271 24052 25283 24055
rect 25774 24052 25780 24064
rect 25271 24024 25780 24052
rect 25271 24021 25283 24024
rect 25225 24015 25283 24021
rect 25774 24012 25780 24024
rect 25832 24012 25838 24064
rect 25958 24012 25964 24064
rect 26016 24052 26022 24064
rect 26605 24055 26663 24061
rect 26605 24052 26617 24055
rect 26016 24024 26617 24052
rect 26016 24012 26022 24024
rect 26605 24021 26617 24024
rect 26651 24021 26663 24055
rect 28810 24052 28816 24064
rect 28723 24024 28816 24052
rect 26605 24015 26663 24021
rect 28810 24012 28816 24024
rect 28868 24052 28874 24064
rect 29638 24052 29644 24064
rect 28868 24024 29644 24052
rect 28868 24012 28874 24024
rect 29638 24012 29644 24024
rect 29696 24012 29702 24064
rect 31202 24012 31208 24064
rect 31260 24052 31266 24064
rect 31297 24055 31355 24061
rect 31297 24052 31309 24055
rect 31260 24024 31309 24052
rect 31260 24012 31266 24024
rect 31297 24021 31309 24024
rect 31343 24021 31355 24055
rect 31726 24052 31754 24092
rect 34808 24064 34836 24092
rect 37274 24080 37280 24092
rect 37332 24080 37338 24132
rect 32398 24052 32404 24064
rect 31726 24024 32404 24052
rect 31297 24015 31355 24021
rect 32398 24012 32404 24024
rect 32456 24012 32462 24064
rect 32493 24055 32551 24061
rect 32493 24021 32505 24055
rect 32539 24052 32551 24055
rect 32950 24052 32956 24064
rect 32539 24024 32956 24052
rect 32539 24021 32551 24024
rect 32493 24015 32551 24021
rect 32950 24012 32956 24024
rect 33008 24012 33014 24064
rect 34790 24052 34796 24064
rect 34703 24024 34796 24052
rect 34790 24012 34796 24024
rect 34848 24012 34854 24064
rect 35529 24055 35587 24061
rect 35529 24021 35541 24055
rect 35575 24052 35587 24055
rect 35618 24052 35624 24064
rect 35575 24024 35624 24052
rect 35575 24021 35587 24024
rect 35529 24015 35587 24021
rect 35618 24012 35624 24024
rect 35676 24012 35682 24064
rect 37734 24052 37740 24064
rect 37695 24024 37740 24052
rect 37734 24012 37740 24024
rect 37792 24012 37798 24064
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 11882 23848 11888 23860
rect 11843 23820 11888 23848
rect 11882 23808 11888 23820
rect 11940 23808 11946 23860
rect 14274 23848 14280 23860
rect 14235 23820 14280 23848
rect 14274 23808 14280 23820
rect 14332 23808 14338 23860
rect 15102 23808 15108 23860
rect 15160 23848 15166 23860
rect 15765 23851 15823 23857
rect 15765 23848 15777 23851
rect 15160 23820 15777 23848
rect 15160 23808 15166 23820
rect 15765 23817 15777 23820
rect 15811 23817 15823 23851
rect 15930 23848 15936 23860
rect 15891 23820 15936 23848
rect 15765 23811 15823 23817
rect 15930 23808 15936 23820
rect 15988 23808 15994 23860
rect 17954 23848 17960 23860
rect 17915 23820 17960 23848
rect 17954 23808 17960 23820
rect 18012 23808 18018 23860
rect 21177 23851 21235 23857
rect 21177 23817 21189 23851
rect 21223 23848 21235 23851
rect 21358 23848 21364 23860
rect 21223 23820 21364 23848
rect 21223 23817 21235 23820
rect 21177 23811 21235 23817
rect 21358 23808 21364 23820
rect 21416 23808 21422 23860
rect 22097 23851 22155 23857
rect 22097 23817 22109 23851
rect 22143 23848 22155 23851
rect 22554 23848 22560 23860
rect 22143 23820 22560 23848
rect 22143 23817 22155 23820
rect 22097 23811 22155 23817
rect 22554 23808 22560 23820
rect 22612 23808 22618 23860
rect 22741 23851 22799 23857
rect 22741 23817 22753 23851
rect 22787 23848 22799 23851
rect 23842 23848 23848 23860
rect 22787 23820 23848 23848
rect 22787 23817 22799 23820
rect 22741 23811 22799 23817
rect 23842 23808 23848 23820
rect 23900 23808 23906 23860
rect 24397 23851 24455 23857
rect 24397 23817 24409 23851
rect 24443 23848 24455 23851
rect 24854 23848 24860 23860
rect 24443 23820 24860 23848
rect 24443 23817 24455 23820
rect 24397 23811 24455 23817
rect 24854 23808 24860 23820
rect 24912 23808 24918 23860
rect 28074 23808 28080 23860
rect 28132 23848 28138 23860
rect 28905 23851 28963 23857
rect 28905 23848 28917 23851
rect 28132 23820 28917 23848
rect 28132 23808 28138 23820
rect 28905 23817 28917 23820
rect 28951 23817 28963 23851
rect 29086 23848 29092 23860
rect 29047 23820 29092 23848
rect 28905 23811 28963 23817
rect 29086 23808 29092 23820
rect 29144 23808 29150 23860
rect 32306 23808 32312 23860
rect 32364 23848 32370 23860
rect 32493 23851 32551 23857
rect 32493 23848 32505 23851
rect 32364 23820 32505 23848
rect 32364 23808 32370 23820
rect 32493 23817 32505 23820
rect 32539 23848 32551 23851
rect 33686 23848 33692 23860
rect 32539 23820 33692 23848
rect 32539 23817 32551 23820
rect 32493 23811 32551 23817
rect 33686 23808 33692 23820
rect 33744 23808 33750 23860
rect 34885 23851 34943 23857
rect 34885 23817 34897 23851
rect 34931 23848 34943 23851
rect 35342 23848 35348 23860
rect 34931 23820 35348 23848
rect 34931 23817 34943 23820
rect 34885 23811 34943 23817
rect 35342 23808 35348 23820
rect 35400 23808 35406 23860
rect 35710 23808 35716 23860
rect 35768 23848 35774 23860
rect 35805 23851 35863 23857
rect 35805 23848 35817 23851
rect 35768 23820 35817 23848
rect 35768 23808 35774 23820
rect 35805 23817 35817 23820
rect 35851 23848 35863 23851
rect 36449 23851 36507 23857
rect 36449 23848 36461 23851
rect 35851 23820 36461 23848
rect 35851 23817 35863 23820
rect 35805 23811 35863 23817
rect 36449 23817 36461 23820
rect 36495 23817 36507 23851
rect 36449 23811 36507 23817
rect 8570 23780 8576 23792
rect 8483 23752 8576 23780
rect 8570 23740 8576 23752
rect 8628 23780 8634 23792
rect 10318 23780 10324 23792
rect 8628 23752 10324 23780
rect 8628 23740 8634 23752
rect 10318 23740 10324 23752
rect 10376 23740 10382 23792
rect 12253 23783 12311 23789
rect 12253 23749 12265 23783
rect 12299 23780 12311 23783
rect 12710 23780 12716 23792
rect 12299 23752 12716 23780
rect 12299 23749 12311 23752
rect 12253 23743 12311 23749
rect 12710 23740 12716 23752
rect 12768 23740 12774 23792
rect 14550 23740 14556 23792
rect 14608 23780 14614 23792
rect 15565 23783 15623 23789
rect 15565 23780 15577 23783
rect 14608 23752 15577 23780
rect 14608 23740 14614 23752
rect 15565 23749 15577 23752
rect 15611 23780 15623 23783
rect 16853 23783 16911 23789
rect 15611 23752 16804 23780
rect 15611 23749 15623 23752
rect 15565 23743 15623 23749
rect 8386 23712 8392 23724
rect 8347 23684 8392 23712
rect 8386 23672 8392 23684
rect 8444 23672 8450 23724
rect 9214 23712 9220 23724
rect 9175 23684 9220 23712
rect 9214 23672 9220 23684
rect 9272 23672 9278 23724
rect 10137 23715 10195 23721
rect 10137 23681 10149 23715
rect 10183 23712 10195 23715
rect 11146 23712 11152 23724
rect 10183 23684 11152 23712
rect 10183 23681 10195 23684
rect 10137 23675 10195 23681
rect 11146 23672 11152 23684
rect 11204 23672 11210 23724
rect 12066 23712 12072 23724
rect 12027 23684 12072 23712
rect 12066 23672 12072 23684
rect 12124 23672 12130 23724
rect 12345 23715 12403 23721
rect 12345 23681 12357 23715
rect 12391 23681 12403 23715
rect 12345 23675 12403 23681
rect 9306 23644 9312 23656
rect 9267 23616 9312 23644
rect 9306 23604 9312 23616
rect 9364 23604 9370 23656
rect 10226 23604 10232 23656
rect 10284 23644 10290 23656
rect 12360 23644 12388 23675
rect 12526 23672 12532 23724
rect 12584 23712 12590 23724
rect 12805 23715 12863 23721
rect 12805 23712 12817 23715
rect 12584 23684 12817 23712
rect 12584 23672 12590 23684
rect 12805 23681 12817 23684
rect 12851 23681 12863 23715
rect 12989 23715 13047 23721
rect 12989 23712 13001 23715
rect 12805 23675 12863 23681
rect 12912 23684 13001 23712
rect 10284 23616 12388 23644
rect 10284 23604 10290 23616
rect 9585 23579 9643 23585
rect 9585 23545 9597 23579
rect 9631 23576 9643 23579
rect 10502 23576 10508 23588
rect 9631 23548 10508 23576
rect 9631 23545 9643 23548
rect 9585 23539 9643 23545
rect 10502 23536 10508 23548
rect 10560 23536 10566 23588
rect 12342 23536 12348 23588
rect 12400 23576 12406 23588
rect 12912 23576 12940 23684
rect 12989 23681 13001 23684
rect 13035 23681 13047 23715
rect 13446 23712 13452 23724
rect 13407 23684 13452 23712
rect 12989 23675 13047 23681
rect 13446 23672 13452 23684
rect 13504 23672 13510 23724
rect 13630 23712 13636 23724
rect 13591 23684 13636 23712
rect 13630 23672 13636 23684
rect 13688 23672 13694 23724
rect 14458 23712 14464 23724
rect 14419 23684 14464 23712
rect 14458 23672 14464 23684
rect 14516 23672 14522 23724
rect 15105 23715 15163 23721
rect 15105 23681 15117 23715
rect 15151 23712 15163 23715
rect 16390 23712 16396 23724
rect 15151 23684 16396 23712
rect 15151 23681 15163 23684
rect 15105 23675 15163 23681
rect 16390 23672 16396 23684
rect 16448 23672 16454 23724
rect 16669 23715 16727 23721
rect 16669 23681 16681 23715
rect 16715 23681 16727 23715
rect 16776 23712 16804 23752
rect 16853 23749 16865 23783
rect 16899 23780 16911 23783
rect 18690 23780 18696 23792
rect 16899 23752 18696 23780
rect 16899 23749 16911 23752
rect 16853 23743 16911 23749
rect 18690 23740 18696 23752
rect 18748 23740 18754 23792
rect 21928 23752 24256 23780
rect 17773 23715 17831 23721
rect 16776 23684 17724 23712
rect 16669 23675 16727 23681
rect 12400 23548 12940 23576
rect 14921 23579 14979 23585
rect 12400 23536 12406 23548
rect 14921 23545 14933 23579
rect 14967 23576 14979 23579
rect 15194 23576 15200 23588
rect 14967 23548 15200 23576
rect 14967 23545 14979 23548
rect 14921 23539 14979 23545
rect 15194 23536 15200 23548
rect 15252 23576 15258 23588
rect 16684 23576 16712 23675
rect 16850 23604 16856 23656
rect 16908 23644 16914 23656
rect 17589 23647 17647 23653
rect 17589 23644 17601 23647
rect 16908 23616 17601 23644
rect 16908 23604 16914 23616
rect 17589 23613 17601 23616
rect 17635 23613 17647 23647
rect 17696 23644 17724 23684
rect 17773 23681 17785 23715
rect 17819 23712 17831 23715
rect 19153 23715 19211 23721
rect 19153 23712 19165 23715
rect 17819 23684 19165 23712
rect 17819 23681 17831 23684
rect 17773 23675 17831 23681
rect 19153 23681 19165 23684
rect 19199 23712 19211 23715
rect 19426 23712 19432 23724
rect 19199 23684 19432 23712
rect 19199 23681 19211 23684
rect 19153 23675 19211 23681
rect 19426 23672 19432 23684
rect 19484 23712 19490 23724
rect 19981 23715 20039 23721
rect 19981 23712 19993 23715
rect 19484 23684 19993 23712
rect 19484 23672 19490 23684
rect 19981 23681 19993 23684
rect 20027 23681 20039 23715
rect 21082 23712 21088 23724
rect 21043 23684 21088 23712
rect 19981 23675 20039 23681
rect 21082 23672 21088 23684
rect 21140 23672 21146 23724
rect 21928 23721 21956 23752
rect 21269 23715 21327 23721
rect 21269 23681 21281 23715
rect 21315 23681 21327 23715
rect 21269 23675 21327 23681
rect 21913 23715 21971 23721
rect 21913 23681 21925 23715
rect 21959 23681 21971 23715
rect 21913 23675 21971 23681
rect 18598 23644 18604 23656
rect 17696 23616 18604 23644
rect 17589 23607 17647 23613
rect 18598 23604 18604 23616
rect 18656 23604 18662 23656
rect 18966 23644 18972 23656
rect 18879 23616 18972 23644
rect 18966 23604 18972 23616
rect 19024 23604 19030 23656
rect 19797 23647 19855 23653
rect 19797 23613 19809 23647
rect 19843 23644 19855 23647
rect 20438 23644 20444 23656
rect 19843 23616 20444 23644
rect 19843 23613 19855 23616
rect 19797 23607 19855 23613
rect 20438 23604 20444 23616
rect 20496 23604 20502 23656
rect 21284 23644 21312 23675
rect 22094 23672 22100 23724
rect 22152 23712 22158 23724
rect 22557 23715 22615 23721
rect 22152 23684 22197 23712
rect 22152 23672 22158 23684
rect 22557 23681 22569 23715
rect 22603 23681 22615 23715
rect 22738 23712 22744 23724
rect 22699 23684 22744 23712
rect 22557 23675 22615 23681
rect 22112 23644 22140 23672
rect 21284 23616 22140 23644
rect 22462 23604 22468 23656
rect 22520 23644 22526 23656
rect 22572 23644 22600 23675
rect 22738 23672 22744 23684
rect 22796 23672 22802 23724
rect 23385 23715 23443 23721
rect 23385 23681 23397 23715
rect 23431 23712 23443 23715
rect 23474 23712 23480 23724
rect 23431 23684 23480 23712
rect 23431 23681 23443 23684
rect 23385 23675 23443 23681
rect 23474 23672 23480 23684
rect 23532 23672 23538 23724
rect 23750 23712 23756 23724
rect 23584 23684 23756 23712
rect 22520 23616 22600 23644
rect 23293 23647 23351 23653
rect 22520 23604 22526 23616
rect 23293 23613 23305 23647
rect 23339 23644 23351 23647
rect 23584 23644 23612 23684
rect 23750 23672 23756 23684
rect 23808 23672 23814 23724
rect 24228 23721 24256 23752
rect 24946 23740 24952 23792
rect 25004 23780 25010 23792
rect 29638 23780 29644 23792
rect 25004 23752 25636 23780
rect 25004 23740 25010 23752
rect 24213 23715 24271 23721
rect 24213 23681 24225 23715
rect 24259 23681 24271 23715
rect 24213 23675 24271 23681
rect 23339 23616 23612 23644
rect 24228 23644 24256 23675
rect 24394 23672 24400 23724
rect 24452 23712 24458 23724
rect 25608 23721 25636 23752
rect 27908 23752 28856 23780
rect 29599 23752 29644 23780
rect 25409 23715 25467 23721
rect 24452 23684 24497 23712
rect 24452 23672 24458 23684
rect 25409 23681 25421 23715
rect 25455 23681 25467 23715
rect 25409 23675 25467 23681
rect 25593 23715 25651 23721
rect 25593 23681 25605 23715
rect 25639 23681 25651 23715
rect 25593 23675 25651 23681
rect 25314 23644 25320 23656
rect 24228 23616 25320 23644
rect 23339 23613 23351 23616
rect 23293 23607 23351 23613
rect 25314 23604 25320 23616
rect 25372 23604 25378 23656
rect 25424 23644 25452 23675
rect 25682 23672 25688 23724
rect 25740 23712 25746 23724
rect 25869 23715 25927 23721
rect 25740 23684 25785 23712
rect 25740 23672 25746 23684
rect 25869 23681 25881 23715
rect 25915 23712 25927 23715
rect 26786 23712 26792 23724
rect 25915 23684 26792 23712
rect 25915 23681 25927 23684
rect 25869 23675 25927 23681
rect 26786 23672 26792 23684
rect 26844 23672 26850 23724
rect 27246 23712 27252 23724
rect 27207 23684 27252 23712
rect 27246 23672 27252 23684
rect 27304 23672 27310 23724
rect 27430 23712 27436 23724
rect 27391 23684 27436 23712
rect 27430 23672 27436 23684
rect 27488 23672 27494 23724
rect 27908 23721 27936 23752
rect 28828 23721 28856 23752
rect 29638 23740 29644 23752
rect 29696 23740 29702 23792
rect 29822 23780 29828 23792
rect 29783 23752 29828 23780
rect 29822 23740 29828 23752
rect 29880 23740 29886 23792
rect 32030 23740 32036 23792
rect 32088 23780 32094 23792
rect 32088 23752 34560 23780
rect 32088 23740 32094 23752
rect 27893 23715 27951 23721
rect 27893 23681 27905 23715
rect 27939 23681 27951 23715
rect 27893 23675 27951 23681
rect 28077 23715 28135 23721
rect 28077 23681 28089 23715
rect 28123 23712 28135 23715
rect 28721 23715 28779 23721
rect 28721 23712 28733 23715
rect 28123 23684 28733 23712
rect 28123 23681 28135 23684
rect 28077 23675 28135 23681
rect 28721 23681 28733 23684
rect 28767 23681 28779 23715
rect 28721 23675 28779 23681
rect 28813 23715 28871 23721
rect 28813 23681 28825 23715
rect 28859 23712 28871 23715
rect 29270 23712 29276 23724
rect 28859 23684 29276 23712
rect 28859 23681 28871 23684
rect 28813 23675 28871 23681
rect 27264 23644 27292 23672
rect 25424 23616 27292 23644
rect 28736 23644 28764 23675
rect 29270 23672 29276 23684
rect 29328 23672 29334 23724
rect 30742 23672 30748 23724
rect 30800 23712 30806 23724
rect 32401 23715 32459 23721
rect 32401 23712 32413 23715
rect 30800 23684 32413 23712
rect 30800 23672 30806 23684
rect 32401 23681 32413 23684
rect 32447 23681 32459 23715
rect 32401 23675 32459 23681
rect 32585 23715 32643 23721
rect 32585 23681 32597 23715
rect 32631 23712 32643 23715
rect 32674 23712 32680 23724
rect 32631 23684 32680 23712
rect 32631 23681 32643 23684
rect 32585 23675 32643 23681
rect 32674 23672 32680 23684
rect 32732 23672 32738 23724
rect 33042 23712 33048 23724
rect 33003 23684 33048 23712
rect 33042 23672 33048 23684
rect 33100 23672 33106 23724
rect 33229 23715 33287 23721
rect 33229 23681 33241 23715
rect 33275 23712 33287 23715
rect 33594 23712 33600 23724
rect 33275 23684 33600 23712
rect 33275 23681 33287 23684
rect 33229 23675 33287 23681
rect 33594 23672 33600 23684
rect 33652 23672 33658 23724
rect 34532 23721 34560 23752
rect 35894 23740 35900 23792
rect 35952 23780 35958 23792
rect 36265 23783 36323 23789
rect 36265 23780 36277 23783
rect 35952 23752 36277 23780
rect 35952 23740 35958 23752
rect 36265 23749 36277 23752
rect 36311 23780 36323 23783
rect 36630 23780 36636 23792
rect 36311 23752 36636 23780
rect 36311 23749 36323 23752
rect 36265 23743 36323 23749
rect 36630 23740 36636 23752
rect 36688 23740 36694 23792
rect 34517 23715 34575 23721
rect 34517 23681 34529 23715
rect 34563 23681 34575 23715
rect 35345 23715 35403 23721
rect 35345 23712 35357 23715
rect 34517 23675 34575 23681
rect 34624 23684 35357 23712
rect 29638 23644 29644 23656
rect 28736 23616 29644 23644
rect 29638 23604 29644 23616
rect 29696 23604 29702 23656
rect 30650 23644 30656 23656
rect 30611 23616 30656 23644
rect 30650 23604 30656 23616
rect 30708 23604 30714 23656
rect 30929 23647 30987 23653
rect 30929 23613 30941 23647
rect 30975 23644 30987 23647
rect 33134 23644 33140 23656
rect 30975 23616 33140 23644
rect 30975 23613 30987 23616
rect 30929 23607 30987 23613
rect 33134 23604 33140 23616
rect 33192 23604 33198 23656
rect 15252 23548 16712 23576
rect 18984 23576 19012 23604
rect 19978 23576 19984 23588
rect 18984 23548 19984 23576
rect 15252 23536 15258 23548
rect 19978 23536 19984 23548
rect 20036 23536 20042 23588
rect 20165 23579 20223 23585
rect 20165 23545 20177 23579
rect 20211 23576 20223 23579
rect 23014 23576 23020 23588
rect 20211 23548 23020 23576
rect 20211 23545 20223 23548
rect 20165 23539 20223 23545
rect 23014 23536 23020 23548
rect 23072 23536 23078 23588
rect 23753 23579 23811 23585
rect 23753 23545 23765 23579
rect 23799 23576 23811 23579
rect 24946 23576 24952 23588
rect 23799 23548 24952 23576
rect 23799 23545 23811 23548
rect 23753 23539 23811 23545
rect 24946 23536 24952 23548
rect 25004 23536 25010 23588
rect 25501 23579 25559 23585
rect 25501 23545 25513 23579
rect 25547 23576 25559 23579
rect 26234 23576 26240 23588
rect 25547 23548 26240 23576
rect 25547 23545 25559 23548
rect 25501 23539 25559 23545
rect 26234 23536 26240 23548
rect 26292 23536 26298 23588
rect 26970 23536 26976 23588
rect 27028 23576 27034 23588
rect 27430 23576 27436 23588
rect 27028 23548 27436 23576
rect 27028 23536 27034 23548
rect 27430 23536 27436 23548
rect 27488 23536 27494 23588
rect 28537 23579 28595 23585
rect 28537 23545 28549 23579
rect 28583 23545 28595 23579
rect 28537 23539 28595 23545
rect 9674 23468 9680 23520
rect 9732 23508 9738 23520
rect 10226 23508 10232 23520
rect 9732 23480 10232 23508
rect 9732 23468 9738 23480
rect 10226 23468 10232 23480
rect 10284 23468 10290 23520
rect 12802 23508 12808 23520
rect 12763 23480 12808 23508
rect 12802 23468 12808 23480
rect 12860 23468 12866 23520
rect 13078 23468 13084 23520
rect 13136 23508 13142 23520
rect 13541 23511 13599 23517
rect 13541 23508 13553 23511
rect 13136 23480 13553 23508
rect 13136 23468 13142 23480
rect 13541 23477 13553 23480
rect 13587 23477 13599 23511
rect 13541 23471 13599 23477
rect 15749 23511 15807 23517
rect 15749 23477 15761 23511
rect 15795 23508 15807 23511
rect 16482 23508 16488 23520
rect 15795 23480 16488 23508
rect 15795 23477 15807 23480
rect 15749 23471 15807 23477
rect 16482 23468 16488 23480
rect 16540 23468 16546 23520
rect 17037 23511 17095 23517
rect 17037 23477 17049 23511
rect 17083 23508 17095 23511
rect 17586 23508 17592 23520
rect 17083 23480 17592 23508
rect 17083 23477 17095 23480
rect 17037 23471 17095 23477
rect 17586 23468 17592 23480
rect 17644 23468 17650 23520
rect 19334 23508 19340 23520
rect 19295 23480 19340 23508
rect 19334 23468 19340 23480
rect 19392 23468 19398 23520
rect 25225 23511 25283 23517
rect 25225 23477 25237 23511
rect 25271 23508 25283 23511
rect 26418 23508 26424 23520
rect 25271 23480 26424 23508
rect 25271 23477 25283 23480
rect 25225 23471 25283 23477
rect 26418 23468 26424 23480
rect 26476 23468 26482 23520
rect 27154 23468 27160 23520
rect 27212 23508 27218 23520
rect 27341 23511 27399 23517
rect 27341 23508 27353 23511
rect 27212 23480 27353 23508
rect 27212 23468 27218 23480
rect 27341 23477 27353 23480
rect 27387 23477 27399 23511
rect 27982 23508 27988 23520
rect 27943 23480 27988 23508
rect 27341 23471 27399 23477
rect 27982 23468 27988 23480
rect 28040 23468 28046 23520
rect 28552 23508 28580 23539
rect 28994 23508 29000 23520
rect 28552 23480 29000 23508
rect 28994 23468 29000 23480
rect 29052 23468 29058 23520
rect 33134 23508 33140 23520
rect 33095 23480 33140 23508
rect 33134 23468 33140 23480
rect 33192 23468 33198 23520
rect 34532 23508 34560 23675
rect 34624 23656 34652 23684
rect 35345 23681 35357 23684
rect 35391 23681 35403 23715
rect 35345 23675 35403 23681
rect 36541 23715 36599 23721
rect 36541 23681 36553 23715
rect 36587 23681 36599 23715
rect 36541 23675 36599 23681
rect 34606 23604 34612 23656
rect 34664 23644 34670 23656
rect 34664 23616 34709 23644
rect 34664 23604 34670 23616
rect 35618 23604 35624 23656
rect 35676 23644 35682 23656
rect 36556 23644 36584 23675
rect 37182 23672 37188 23724
rect 37240 23712 37246 23724
rect 37461 23715 37519 23721
rect 37461 23712 37473 23715
rect 37240 23684 37473 23712
rect 37240 23672 37246 23684
rect 37461 23681 37473 23684
rect 37507 23681 37519 23715
rect 37461 23675 37519 23681
rect 35676 23616 36584 23644
rect 37553 23647 37611 23653
rect 35676 23604 35682 23616
rect 37553 23613 37565 23647
rect 37599 23644 37611 23647
rect 37734 23644 37740 23656
rect 37599 23616 37740 23644
rect 37599 23613 37611 23616
rect 37553 23607 37611 23613
rect 37734 23604 37740 23616
rect 37792 23604 37798 23656
rect 35437 23511 35495 23517
rect 35437 23508 35449 23511
rect 34532 23480 35449 23508
rect 35437 23477 35449 23480
rect 35483 23477 35495 23511
rect 35437 23471 35495 23477
rect 36265 23511 36323 23517
rect 36265 23477 36277 23511
rect 36311 23508 36323 23511
rect 36722 23508 36728 23520
rect 36311 23480 36728 23508
rect 36311 23477 36323 23480
rect 36265 23471 36323 23477
rect 36722 23468 36728 23480
rect 36780 23468 36786 23520
rect 37826 23508 37832 23520
rect 37787 23480 37832 23508
rect 37826 23468 37832 23480
rect 37884 23468 37890 23520
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 8386 23304 8392 23316
rect 8347 23276 8392 23304
rect 8386 23264 8392 23276
rect 8444 23264 8450 23316
rect 9214 23264 9220 23316
rect 9272 23304 9278 23316
rect 9493 23307 9551 23313
rect 9493 23304 9505 23307
rect 9272 23276 9505 23304
rect 9272 23264 9278 23276
rect 9493 23273 9505 23276
rect 9539 23273 9551 23307
rect 9493 23267 9551 23273
rect 11609 23307 11667 23313
rect 11609 23273 11621 23307
rect 11655 23304 11667 23307
rect 12526 23304 12532 23316
rect 11655 23276 12532 23304
rect 11655 23273 11667 23276
rect 11609 23267 11667 23273
rect 12526 23264 12532 23276
rect 12584 23264 12590 23316
rect 15010 23264 15016 23316
rect 15068 23304 15074 23316
rect 18782 23304 18788 23316
rect 15068 23276 18788 23304
rect 15068 23264 15074 23276
rect 18782 23264 18788 23276
rect 18840 23264 18846 23316
rect 20990 23304 20996 23316
rect 20456 23276 20996 23304
rect 10594 23196 10600 23248
rect 10652 23236 10658 23248
rect 12250 23236 12256 23248
rect 10652 23208 12256 23236
rect 10652 23196 10658 23208
rect 12250 23196 12256 23208
rect 12308 23236 12314 23248
rect 12308 23208 13124 23236
rect 12308 23196 12314 23208
rect 9030 23128 9036 23180
rect 9088 23168 9094 23180
rect 9217 23171 9275 23177
rect 9217 23168 9229 23171
rect 9088 23140 9229 23168
rect 9088 23128 9094 23140
rect 9217 23137 9229 23140
rect 9263 23168 9275 23171
rect 11146 23168 11152 23180
rect 9263 23140 11152 23168
rect 9263 23137 9275 23140
rect 9217 23131 9275 23137
rect 11146 23128 11152 23140
rect 11204 23128 11210 23180
rect 11974 23128 11980 23180
rect 12032 23168 12038 23180
rect 12032 23140 12848 23168
rect 12032 23128 12038 23140
rect 7006 23100 7012 23112
rect 6967 23072 7012 23100
rect 7006 23060 7012 23072
rect 7064 23060 7070 23112
rect 8386 23060 8392 23112
rect 8444 23100 8450 23112
rect 8938 23100 8944 23112
rect 8444 23072 8944 23100
rect 8444 23060 8450 23072
rect 8938 23060 8944 23072
rect 8996 23100 9002 23112
rect 9125 23103 9183 23109
rect 9125 23100 9137 23103
rect 8996 23072 9137 23100
rect 8996 23060 9002 23072
rect 9125 23069 9137 23072
rect 9171 23069 9183 23103
rect 10226 23100 10232 23112
rect 10187 23072 10232 23100
rect 9125 23063 9183 23069
rect 10226 23060 10232 23072
rect 10284 23060 10290 23112
rect 10321 23103 10379 23109
rect 10321 23069 10333 23103
rect 10367 23069 10379 23103
rect 10321 23063 10379 23069
rect 7276 23035 7334 23041
rect 7276 23001 7288 23035
rect 7322 23032 7334 23035
rect 9953 23035 10011 23041
rect 9953 23032 9965 23035
rect 7322 23004 9965 23032
rect 7322 23001 7334 23004
rect 7276 22995 7334 23001
rect 9953 23001 9965 23004
rect 9999 23001 10011 23035
rect 9953 22995 10011 23001
rect 10336 22964 10364 23063
rect 10410 23060 10416 23112
rect 10468 23100 10474 23112
rect 10468 23072 10513 23100
rect 10468 23060 10474 23072
rect 10594 23060 10600 23112
rect 10652 23100 10658 23112
rect 11241 23103 11299 23109
rect 10652 23072 10697 23100
rect 10652 23060 10658 23072
rect 11241 23069 11253 23103
rect 11287 23100 11299 23103
rect 12710 23100 12716 23112
rect 11287 23072 12204 23100
rect 12671 23072 12716 23100
rect 11287 23069 11299 23072
rect 11241 23063 11299 23069
rect 11054 22964 11060 22976
rect 10336 22936 11060 22964
rect 11054 22924 11060 22936
rect 11112 22924 11118 22976
rect 12176 22964 12204 23072
rect 12710 23060 12716 23072
rect 12768 23060 12774 23112
rect 12820 23109 12848 23140
rect 12805 23103 12863 23109
rect 12805 23069 12817 23103
rect 12851 23069 12863 23103
rect 12805 23063 12863 23069
rect 12894 23060 12900 23112
rect 12952 23100 12958 23112
rect 13096 23109 13124 23208
rect 15102 23196 15108 23248
rect 15160 23236 15166 23248
rect 17770 23236 17776 23248
rect 15160 23208 17080 23236
rect 17731 23208 17776 23236
rect 15160 23196 15166 23208
rect 13081 23103 13139 23109
rect 12952 23072 12997 23100
rect 12952 23060 12958 23072
rect 13081 23069 13093 23103
rect 13127 23069 13139 23103
rect 13081 23063 13139 23069
rect 13170 23060 13176 23112
rect 13228 23100 13234 23112
rect 14093 23103 14151 23109
rect 14093 23100 14105 23103
rect 13228 23072 14105 23100
rect 13228 23060 13234 23072
rect 14093 23069 14105 23072
rect 14139 23069 14151 23103
rect 16758 23100 16764 23112
rect 16719 23072 16764 23100
rect 14093 23063 14151 23069
rect 16758 23060 16764 23072
rect 16816 23060 16822 23112
rect 17052 23109 17080 23208
rect 17770 23196 17776 23208
rect 17828 23196 17834 23248
rect 19613 23171 19671 23177
rect 19613 23168 19625 23171
rect 18708 23140 19625 23168
rect 17037 23103 17095 23109
rect 17037 23069 17049 23103
rect 17083 23069 17095 23103
rect 17586 23100 17592 23112
rect 17547 23072 17592 23100
rect 17037 23063 17095 23069
rect 17586 23060 17592 23072
rect 17644 23060 17650 23112
rect 18708 23109 18736 23140
rect 19613 23137 19625 23140
rect 19659 23137 19671 23171
rect 19613 23131 19671 23137
rect 20254 23128 20260 23180
rect 20312 23168 20318 23180
rect 20456 23177 20484 23276
rect 20990 23264 20996 23276
rect 21048 23264 21054 23316
rect 26053 23307 26111 23313
rect 26053 23273 26065 23307
rect 26099 23304 26111 23307
rect 26602 23304 26608 23316
rect 26099 23276 26608 23304
rect 26099 23273 26111 23276
rect 26053 23267 26111 23273
rect 26602 23264 26608 23276
rect 26660 23264 26666 23316
rect 26786 23304 26792 23316
rect 26747 23276 26792 23304
rect 26786 23264 26792 23276
rect 26844 23264 26850 23316
rect 27798 23264 27804 23316
rect 27856 23304 27862 23316
rect 28534 23304 28540 23316
rect 27856 23276 28540 23304
rect 27856 23264 27862 23276
rect 28534 23264 28540 23276
rect 28592 23264 28598 23316
rect 31478 23304 31484 23316
rect 30484 23276 31156 23304
rect 31439 23276 31484 23304
rect 21008 23236 21036 23264
rect 21726 23236 21732 23248
rect 21008 23208 21732 23236
rect 21726 23196 21732 23208
rect 21784 23236 21790 23248
rect 24670 23236 24676 23248
rect 21784 23208 22048 23236
rect 21784 23196 21790 23208
rect 22020 23177 22048 23208
rect 23676 23208 24676 23236
rect 20441 23171 20499 23177
rect 20441 23168 20453 23171
rect 20312 23140 20453 23168
rect 20312 23128 20318 23140
rect 20441 23137 20453 23140
rect 20487 23137 20499 23171
rect 22005 23171 22063 23177
rect 20441 23131 20499 23137
rect 21100 23140 21680 23168
rect 18693 23103 18751 23109
rect 18693 23069 18705 23103
rect 18739 23069 18751 23103
rect 18693 23063 18751 23069
rect 18782 23060 18788 23112
rect 18840 23100 18846 23112
rect 19245 23103 19303 23109
rect 19245 23100 19257 23103
rect 18840 23072 19257 23100
rect 18840 23060 18846 23072
rect 19245 23069 19257 23072
rect 19291 23069 19303 23103
rect 19426 23100 19432 23112
rect 19387 23072 19432 23100
rect 19245 23063 19303 23069
rect 19426 23060 19432 23072
rect 19484 23060 19490 23112
rect 20717 23103 20775 23109
rect 20717 23069 20729 23103
rect 20763 23069 20775 23103
rect 20717 23063 20775 23069
rect 12437 23035 12495 23041
rect 12437 23001 12449 23035
rect 12483 23032 12495 23035
rect 14338 23035 14396 23041
rect 14338 23032 14350 23035
rect 12483 23004 14350 23032
rect 12483 23001 12495 23004
rect 12437 22995 12495 23001
rect 14338 23001 14350 23004
rect 14384 23001 14396 23035
rect 14338 22995 14396 23001
rect 16577 23035 16635 23041
rect 16577 23001 16589 23035
rect 16623 23032 16635 23035
rect 17954 23032 17960 23044
rect 16623 23004 17960 23032
rect 16623 23001 16635 23004
rect 16577 22995 16635 23001
rect 17954 22992 17960 23004
rect 18012 22992 18018 23044
rect 20732 23032 20760 23063
rect 20806 23060 20812 23112
rect 20864 23100 20870 23112
rect 21100 23100 21128 23140
rect 21542 23100 21548 23112
rect 20864 23072 21128 23100
rect 21503 23072 21548 23100
rect 20864 23060 20870 23072
rect 21542 23060 21548 23072
rect 21600 23060 21606 23112
rect 21652 23100 21680 23140
rect 22005 23137 22017 23171
rect 22051 23137 22063 23171
rect 23676 23168 23704 23208
rect 24670 23196 24676 23208
rect 24728 23236 24734 23248
rect 24765 23239 24823 23245
rect 24765 23236 24777 23239
rect 24728 23208 24777 23236
rect 24728 23196 24734 23208
rect 24765 23205 24777 23208
rect 24811 23205 24823 23239
rect 24765 23199 24823 23205
rect 25682 23196 25688 23248
rect 25740 23236 25746 23248
rect 27709 23239 27767 23245
rect 25740 23208 27660 23236
rect 25740 23196 25746 23208
rect 25501 23171 25559 23177
rect 22005 23131 22063 23137
rect 23584 23140 23704 23168
rect 23768 23140 25452 23168
rect 22281 23103 22339 23109
rect 22281 23100 22293 23103
rect 21652 23072 22293 23100
rect 22281 23069 22293 23072
rect 22327 23069 22339 23103
rect 22281 23063 22339 23069
rect 23474 23060 23480 23112
rect 23532 23100 23538 23112
rect 23584 23109 23612 23140
rect 23569 23103 23627 23109
rect 23569 23100 23581 23103
rect 23532 23072 23581 23100
rect 23532 23060 23538 23072
rect 23569 23069 23581 23072
rect 23615 23069 23627 23103
rect 23768 23100 23796 23140
rect 25424 23112 25452 23140
rect 25501 23137 25513 23171
rect 25547 23168 25559 23171
rect 25547 23140 26372 23168
rect 25547 23137 25559 23140
rect 25501 23131 25559 23137
rect 23569 23063 23627 23069
rect 23672 23072 23796 23100
rect 24765 23103 24823 23109
rect 18524 23004 20760 23032
rect 12618 22964 12624 22976
rect 12176 22936 12624 22964
rect 12618 22924 12624 22936
rect 12676 22964 12682 22976
rect 14826 22964 14832 22976
rect 12676 22936 14832 22964
rect 12676 22924 12682 22936
rect 14826 22924 14832 22936
rect 14884 22964 14890 22976
rect 15473 22967 15531 22973
rect 15473 22964 15485 22967
rect 14884 22936 15485 22964
rect 14884 22924 14890 22936
rect 15473 22933 15485 22936
rect 15519 22933 15531 22967
rect 15473 22927 15531 22933
rect 16390 22924 16396 22976
rect 16448 22964 16454 22976
rect 18524 22973 18552 23004
rect 22738 22992 22744 23044
rect 22796 23032 22802 23044
rect 23672 23032 23700 23072
rect 24765 23069 24777 23103
rect 24811 23069 24823 23103
rect 24765 23063 24823 23069
rect 24949 23103 25007 23109
rect 24949 23069 24961 23103
rect 24995 23100 25007 23103
rect 25038 23100 25044 23112
rect 24995 23072 25044 23100
rect 24995 23069 25007 23072
rect 24949 23063 25007 23069
rect 22796 23004 23700 23032
rect 22796 22992 22802 23004
rect 23750 22992 23756 23044
rect 23808 23032 23814 23044
rect 24780 23032 24808 23063
rect 25038 23060 25044 23072
rect 25096 23060 25102 23112
rect 25406 23100 25412 23112
rect 25367 23072 25412 23100
rect 25406 23060 25412 23072
rect 25464 23060 25470 23112
rect 25593 23103 25651 23109
rect 25593 23069 25605 23103
rect 25639 23100 25651 23103
rect 25866 23100 25872 23112
rect 25639 23072 25872 23100
rect 25639 23069 25651 23072
rect 25593 23063 25651 23069
rect 25866 23060 25872 23072
rect 25924 23060 25930 23112
rect 26234 23060 26240 23112
rect 26292 23060 26298 23112
rect 26344 23109 26372 23140
rect 26602 23128 26608 23180
rect 26660 23168 26666 23180
rect 27522 23168 27528 23180
rect 26660 23140 27528 23168
rect 26660 23128 26666 23140
rect 27522 23128 27528 23140
rect 27580 23128 27586 23180
rect 27632 23168 27660 23208
rect 27709 23205 27721 23239
rect 27755 23236 27767 23239
rect 28074 23236 28080 23248
rect 27755 23208 28080 23236
rect 27755 23205 27767 23208
rect 27709 23199 27767 23205
rect 28074 23196 28080 23208
rect 28132 23196 28138 23248
rect 28350 23168 28356 23180
rect 27632 23140 28356 23168
rect 28350 23128 28356 23140
rect 28408 23128 28414 23180
rect 28445 23171 28503 23177
rect 28445 23137 28457 23171
rect 28491 23168 28503 23171
rect 28994 23168 29000 23180
rect 28491 23140 29000 23168
rect 28491 23137 28503 23140
rect 28445 23131 28503 23137
rect 28994 23128 29000 23140
rect 29052 23128 29058 23180
rect 29362 23168 29368 23180
rect 29104 23140 29368 23168
rect 26329 23103 26387 23109
rect 26329 23069 26341 23103
rect 26375 23069 26387 23103
rect 26329 23063 26387 23069
rect 26789 23103 26847 23109
rect 26789 23069 26801 23103
rect 26835 23069 26847 23103
rect 26789 23063 26847 23069
rect 26053 23035 26111 23041
rect 26053 23032 26065 23035
rect 23808 23004 23853 23032
rect 24780 23004 26065 23032
rect 23808 22992 23814 23004
rect 26053 23001 26065 23004
rect 26099 23032 26111 23035
rect 26252 23032 26280 23060
rect 26804 23032 26832 23063
rect 26878 23060 26884 23112
rect 26936 23100 26942 23112
rect 26973 23103 27031 23109
rect 26973 23100 26985 23103
rect 26936 23072 26985 23100
rect 26936 23060 26942 23072
rect 26973 23069 26985 23072
rect 27019 23069 27031 23103
rect 26973 23063 27031 23069
rect 27617 23103 27675 23109
rect 27617 23069 27629 23103
rect 27663 23069 27675 23103
rect 27798 23100 27804 23112
rect 27759 23072 27804 23100
rect 27617 23063 27675 23069
rect 27062 23032 27068 23044
rect 26099 23004 27068 23032
rect 26099 23001 26111 23004
rect 26053 22995 26111 23001
rect 27062 22992 27068 23004
rect 27120 22992 27126 23044
rect 27632 23032 27660 23063
rect 27798 23060 27804 23072
rect 27856 23060 27862 23112
rect 27982 23060 27988 23112
rect 28040 23100 28046 23112
rect 28261 23103 28319 23109
rect 28261 23100 28273 23103
rect 28040 23072 28273 23100
rect 28040 23060 28046 23072
rect 28261 23069 28273 23072
rect 28307 23069 28319 23103
rect 28261 23063 28319 23069
rect 28537 23103 28595 23109
rect 28537 23069 28549 23103
rect 28583 23100 28595 23103
rect 28810 23100 28816 23112
rect 28583 23072 28816 23100
rect 28583 23069 28595 23072
rect 28537 23063 28595 23069
rect 28810 23060 28816 23072
rect 28868 23060 28874 23112
rect 29104 23100 29132 23140
rect 29362 23128 29368 23140
rect 29420 23168 29426 23180
rect 29733 23171 29791 23177
rect 29733 23168 29745 23171
rect 29420 23140 29745 23168
rect 29420 23128 29426 23140
rect 29733 23137 29745 23140
rect 29779 23137 29791 23171
rect 30374 23168 30380 23180
rect 30335 23140 30380 23168
rect 29733 23131 29791 23137
rect 30374 23128 30380 23140
rect 30432 23128 30438 23180
rect 30484 23109 30512 23276
rect 30837 23239 30895 23245
rect 30837 23205 30849 23239
rect 30883 23205 30895 23239
rect 31128 23236 31156 23276
rect 31478 23264 31484 23276
rect 31536 23264 31542 23316
rect 31849 23307 31907 23313
rect 31849 23273 31861 23307
rect 31895 23304 31907 23307
rect 33042 23304 33048 23316
rect 31895 23276 33048 23304
rect 31895 23273 31907 23276
rect 31849 23267 31907 23273
rect 33042 23264 33048 23276
rect 33100 23264 33106 23316
rect 35618 23264 35624 23316
rect 35676 23304 35682 23316
rect 35897 23307 35955 23313
rect 35897 23304 35909 23307
rect 35676 23276 35909 23304
rect 35676 23264 35682 23276
rect 35897 23273 35909 23276
rect 35943 23273 35955 23307
rect 36722 23304 36728 23316
rect 36683 23276 36728 23304
rect 35897 23267 35955 23273
rect 36722 23264 36728 23276
rect 36780 23264 36786 23316
rect 37090 23304 37096 23316
rect 37051 23276 37096 23304
rect 37090 23264 37096 23276
rect 37148 23264 37154 23316
rect 37642 23304 37648 23316
rect 37603 23276 37648 23304
rect 37642 23264 37648 23276
rect 37700 23264 37706 23316
rect 32122 23236 32128 23248
rect 31128 23208 32128 23236
rect 30837 23199 30895 23205
rect 28920 23072 29132 23100
rect 29641 23103 29699 23109
rect 28626 23032 28632 23044
rect 27632 23004 28632 23032
rect 28626 22992 28632 23004
rect 28684 23032 28690 23044
rect 28920 23032 28948 23072
rect 29641 23069 29653 23103
rect 29687 23069 29699 23103
rect 29641 23063 29699 23069
rect 29825 23103 29883 23109
rect 29825 23069 29837 23103
rect 29871 23069 29883 23103
rect 29825 23063 29883 23069
rect 30469 23103 30527 23109
rect 30469 23069 30481 23103
rect 30515 23069 30527 23103
rect 30852 23100 30880 23199
rect 32122 23196 32128 23208
rect 32180 23196 32186 23248
rect 31573 23171 31631 23177
rect 31573 23137 31585 23171
rect 31619 23168 31631 23171
rect 31938 23168 31944 23180
rect 31619 23140 31944 23168
rect 31619 23137 31631 23140
rect 31573 23131 31631 23137
rect 31938 23128 31944 23140
rect 31996 23128 32002 23180
rect 31478 23100 31484 23112
rect 30852 23072 31484 23100
rect 30469 23063 30527 23069
rect 28684 23004 28948 23032
rect 28684 22992 28690 23004
rect 16945 22967 17003 22973
rect 16945 22964 16957 22967
rect 16448 22936 16957 22964
rect 16448 22924 16454 22936
rect 16945 22933 16957 22936
rect 16991 22933 17003 22967
rect 16945 22927 17003 22933
rect 18509 22967 18567 22973
rect 18509 22933 18521 22967
rect 18555 22933 18567 22967
rect 18509 22927 18567 22933
rect 23017 22967 23075 22973
rect 23017 22933 23029 22967
rect 23063 22964 23075 22967
rect 25682 22964 25688 22976
rect 23063 22936 25688 22964
rect 23063 22933 23075 22936
rect 23017 22927 23075 22933
rect 25682 22924 25688 22936
rect 25740 22924 25746 22976
rect 26237 22967 26295 22973
rect 26237 22933 26249 22967
rect 26283 22964 26295 22967
rect 26326 22964 26332 22976
rect 26283 22936 26332 22964
rect 26283 22933 26295 22936
rect 26237 22927 26295 22933
rect 26326 22924 26332 22936
rect 26384 22924 26390 22976
rect 27246 22924 27252 22976
rect 27304 22964 27310 22976
rect 28721 22967 28779 22973
rect 28721 22964 28733 22967
rect 27304 22936 28733 22964
rect 27304 22924 27310 22936
rect 28721 22933 28733 22936
rect 28767 22933 28779 22967
rect 29656 22964 29684 23063
rect 29840 23032 29868 23063
rect 31478 23060 31484 23072
rect 31536 23060 31542 23112
rect 32769 23103 32827 23109
rect 32769 23069 32781 23103
rect 32815 23100 32827 23103
rect 33134 23100 33140 23112
rect 32815 23072 33140 23100
rect 32815 23069 32827 23072
rect 32769 23063 32827 23069
rect 33134 23060 33140 23072
rect 33192 23060 33198 23112
rect 33686 23100 33692 23112
rect 33647 23072 33692 23100
rect 33686 23060 33692 23072
rect 33744 23060 33750 23112
rect 34885 23103 34943 23109
rect 34885 23069 34897 23103
rect 34931 23100 34943 23103
rect 35342 23100 35348 23112
rect 34931 23072 35348 23100
rect 34931 23069 34943 23072
rect 34885 23063 34943 23069
rect 35342 23060 35348 23072
rect 35400 23060 35406 23112
rect 36630 23100 36636 23112
rect 36591 23072 36636 23100
rect 36630 23060 36636 23072
rect 36688 23060 36694 23112
rect 37553 23103 37611 23109
rect 37553 23069 37565 23103
rect 37599 23100 37611 23103
rect 37734 23100 37740 23112
rect 37599 23072 37740 23100
rect 37599 23069 37611 23072
rect 37553 23063 37611 23069
rect 37734 23060 37740 23072
rect 37792 23060 37798 23112
rect 30834 23032 30840 23044
rect 29840 23004 30840 23032
rect 30834 22992 30840 23004
rect 30892 22992 30898 23044
rect 32950 23032 32956 23044
rect 32911 23004 32956 23032
rect 32950 22992 32956 23004
rect 33008 22992 33014 23044
rect 34790 22992 34796 23044
rect 34848 23032 34854 23044
rect 35069 23035 35127 23041
rect 35069 23032 35081 23035
rect 34848 23004 35081 23032
rect 34848 22992 34854 23004
rect 35069 23001 35081 23004
rect 35115 23001 35127 23035
rect 35710 23032 35716 23044
rect 35671 23004 35716 23032
rect 35069 22995 35127 23001
rect 35710 22992 35716 23004
rect 35768 22992 35774 23044
rect 31018 22964 31024 22976
rect 29656 22936 31024 22964
rect 28721 22927 28779 22933
rect 31018 22924 31024 22936
rect 31076 22924 31082 22976
rect 33137 22967 33195 22973
rect 33137 22933 33149 22967
rect 33183 22964 33195 22967
rect 33226 22964 33232 22976
rect 33183 22936 33232 22964
rect 33183 22933 33195 22936
rect 33137 22927 33195 22933
rect 33226 22924 33232 22936
rect 33284 22924 33290 22976
rect 33410 22924 33416 22976
rect 33468 22964 33474 22976
rect 33778 22964 33784 22976
rect 33468 22936 33784 22964
rect 33468 22924 33474 22936
rect 33778 22924 33784 22936
rect 33836 22924 33842 22976
rect 35253 22967 35311 22973
rect 35253 22933 35265 22967
rect 35299 22964 35311 22967
rect 35434 22964 35440 22976
rect 35299 22936 35440 22964
rect 35299 22933 35311 22936
rect 35253 22927 35311 22933
rect 35434 22924 35440 22936
rect 35492 22924 35498 22976
rect 35894 22924 35900 22976
rect 35952 22973 35958 22976
rect 35952 22967 35971 22973
rect 35959 22933 35971 22967
rect 36078 22964 36084 22976
rect 36039 22936 36084 22964
rect 35952 22927 35971 22933
rect 35952 22924 35958 22927
rect 36078 22924 36084 22936
rect 36136 22924 36142 22976
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 9306 22720 9312 22772
rect 9364 22760 9370 22772
rect 9585 22763 9643 22769
rect 9585 22760 9597 22763
rect 9364 22732 9597 22760
rect 9364 22720 9370 22732
rect 9585 22729 9597 22732
rect 9631 22729 9643 22763
rect 9585 22723 9643 22729
rect 10410 22720 10416 22772
rect 10468 22760 10474 22772
rect 10597 22763 10655 22769
rect 10597 22760 10609 22763
rect 10468 22732 10609 22760
rect 10468 22720 10474 22732
rect 10597 22729 10609 22732
rect 10643 22729 10655 22763
rect 10597 22723 10655 22729
rect 12066 22720 12072 22772
rect 12124 22760 12130 22772
rect 12345 22763 12403 22769
rect 12345 22760 12357 22763
rect 12124 22732 12357 22760
rect 12124 22720 12130 22732
rect 12345 22729 12357 22732
rect 12391 22729 12403 22763
rect 12345 22723 12403 22729
rect 12360 22692 12388 22723
rect 12894 22720 12900 22772
rect 12952 22760 12958 22772
rect 13081 22763 13139 22769
rect 13081 22760 13093 22763
rect 12952 22732 13093 22760
rect 12952 22720 12958 22732
rect 13081 22729 13093 22732
rect 13127 22729 13139 22763
rect 13081 22723 13139 22729
rect 16758 22720 16764 22772
rect 16816 22760 16822 22772
rect 17589 22763 17647 22769
rect 17589 22760 17601 22763
rect 16816 22732 17601 22760
rect 16816 22720 16822 22732
rect 17589 22729 17601 22732
rect 17635 22760 17647 22763
rect 17678 22760 17684 22772
rect 17635 22732 17684 22760
rect 17635 22729 17647 22732
rect 17589 22723 17647 22729
rect 17678 22720 17684 22732
rect 17736 22760 17742 22772
rect 19426 22760 19432 22772
rect 17736 22732 19432 22760
rect 17736 22720 17742 22732
rect 14274 22692 14280 22704
rect 8772 22664 9812 22692
rect 12360 22664 12940 22692
rect 14187 22664 14280 22692
rect 8772 22633 8800 22664
rect 8757 22627 8815 22633
rect 8757 22593 8769 22627
rect 8803 22593 8815 22627
rect 8938 22624 8944 22636
rect 8899 22596 8944 22624
rect 8757 22587 8815 22593
rect 8938 22584 8944 22596
rect 8996 22584 9002 22636
rect 9030 22584 9036 22636
rect 9088 22624 9094 22636
rect 9784 22633 9812 22664
rect 9769 22627 9827 22633
rect 9088 22596 9133 22624
rect 9088 22584 9094 22596
rect 9769 22593 9781 22627
rect 9815 22624 9827 22627
rect 9858 22624 9864 22636
rect 9815 22596 9864 22624
rect 9815 22593 9827 22596
rect 9769 22587 9827 22593
rect 9858 22584 9864 22596
rect 9916 22584 9922 22636
rect 10042 22624 10048 22636
rect 10003 22596 10048 22624
rect 10042 22584 10048 22596
rect 10100 22584 10106 22636
rect 10502 22624 10508 22636
rect 10463 22596 10508 22624
rect 10502 22584 10508 22596
rect 10560 22584 10566 22636
rect 10689 22627 10747 22633
rect 10689 22593 10701 22627
rect 10735 22624 10747 22627
rect 11054 22624 11060 22636
rect 10735 22596 11060 22624
rect 10735 22593 10747 22596
rect 10689 22587 10747 22593
rect 11054 22584 11060 22596
rect 11112 22624 11118 22636
rect 12066 22624 12072 22636
rect 11112 22596 12072 22624
rect 11112 22584 11118 22596
rect 12066 22584 12072 22596
rect 12124 22584 12130 22636
rect 12161 22627 12219 22633
rect 12161 22593 12173 22627
rect 12207 22624 12219 22627
rect 12434 22624 12440 22636
rect 12207 22596 12440 22624
rect 12207 22593 12219 22596
rect 12161 22587 12219 22593
rect 12434 22584 12440 22596
rect 12492 22584 12498 22636
rect 12802 22624 12808 22636
rect 12763 22596 12808 22624
rect 12802 22584 12808 22596
rect 12860 22584 12866 22636
rect 12912 22633 12940 22664
rect 14274 22652 14280 22664
rect 14332 22692 14338 22704
rect 14550 22692 14556 22704
rect 14332 22664 14556 22692
rect 14332 22652 14338 22664
rect 14550 22652 14556 22664
rect 14608 22652 14614 22704
rect 14826 22692 14832 22704
rect 14787 22664 14832 22692
rect 14826 22652 14832 22664
rect 14884 22652 14890 22704
rect 16669 22695 16727 22701
rect 16669 22661 16681 22695
rect 16715 22692 16727 22695
rect 18506 22692 18512 22704
rect 16715 22664 18512 22692
rect 16715 22661 16727 22664
rect 16669 22655 16727 22661
rect 12897 22627 12955 22633
rect 12897 22593 12909 22627
rect 12943 22593 12955 22627
rect 14093 22627 14151 22633
rect 12897 22587 12955 22593
rect 13004 22596 13768 22624
rect 8846 22516 8852 22568
rect 8904 22556 8910 22568
rect 11977 22559 12035 22565
rect 8904 22528 8949 22556
rect 8904 22516 8910 22528
rect 11977 22525 11989 22559
rect 12023 22556 12035 22559
rect 12342 22556 12348 22568
rect 12023 22528 12348 22556
rect 12023 22525 12035 22528
rect 11977 22519 12035 22525
rect 12342 22516 12348 22528
rect 12400 22516 12406 22568
rect 12710 22516 12716 22568
rect 12768 22556 12774 22568
rect 13004 22556 13032 22596
rect 12768 22528 13032 22556
rect 13081 22559 13139 22565
rect 12768 22516 12774 22528
rect 13081 22525 13093 22559
rect 13127 22556 13139 22559
rect 13630 22556 13636 22568
rect 13127 22528 13636 22556
rect 13127 22525 13139 22528
rect 13081 22519 13139 22525
rect 8573 22423 8631 22429
rect 8573 22389 8585 22423
rect 8619 22420 8631 22423
rect 8754 22420 8760 22432
rect 8619 22392 8760 22420
rect 8619 22389 8631 22392
rect 8573 22383 8631 22389
rect 8754 22380 8760 22392
rect 8812 22380 8818 22432
rect 9674 22380 9680 22432
rect 9732 22420 9738 22432
rect 9953 22423 10011 22429
rect 9953 22420 9965 22423
rect 9732 22392 9965 22420
rect 9732 22380 9738 22392
rect 9953 22389 9965 22392
rect 9999 22389 10011 22423
rect 9953 22383 10011 22389
rect 12066 22380 12072 22432
rect 12124 22420 12130 22432
rect 13096 22420 13124 22519
rect 13630 22516 13636 22528
rect 13688 22516 13694 22568
rect 13740 22556 13768 22596
rect 14093 22593 14105 22627
rect 14139 22624 14151 22627
rect 14366 22624 14372 22636
rect 14139 22596 14372 22624
rect 14139 22593 14151 22596
rect 14093 22587 14151 22593
rect 14366 22584 14372 22596
rect 14424 22584 14430 22636
rect 15470 22584 15476 22636
rect 15528 22624 15534 22636
rect 15565 22627 15623 22633
rect 15565 22624 15577 22627
rect 15528 22596 15577 22624
rect 15528 22584 15534 22596
rect 15565 22593 15577 22596
rect 15611 22593 15623 22627
rect 15565 22587 15623 22593
rect 16390 22584 16396 22636
rect 16448 22624 16454 22636
rect 17788 22633 17816 22664
rect 18506 22652 18512 22664
rect 18564 22652 18570 22704
rect 16853 22627 16911 22633
rect 16853 22624 16865 22627
rect 16448 22596 16865 22624
rect 16448 22584 16454 22596
rect 16853 22593 16865 22596
rect 16899 22624 16911 22627
rect 17773 22627 17831 22633
rect 16899 22596 17724 22624
rect 16899 22593 16911 22596
rect 16853 22587 16911 22593
rect 15013 22559 15071 22565
rect 15013 22556 15025 22559
rect 13740 22528 15025 22556
rect 15013 22525 15025 22528
rect 15059 22556 15071 22559
rect 15654 22556 15660 22568
rect 15059 22528 15660 22556
rect 15059 22525 15071 22528
rect 15013 22519 15071 22525
rect 15654 22516 15660 22528
rect 15712 22516 15718 22568
rect 16945 22559 17003 22565
rect 16945 22525 16957 22559
rect 16991 22525 17003 22559
rect 16945 22519 17003 22525
rect 15286 22448 15292 22500
rect 15344 22488 15350 22500
rect 16960 22488 16988 22519
rect 17034 22516 17040 22568
rect 17092 22556 17098 22568
rect 17696 22556 17724 22596
rect 17773 22593 17785 22627
rect 17819 22593 17831 22627
rect 17773 22587 17831 22593
rect 18417 22627 18475 22633
rect 18417 22593 18429 22627
rect 18463 22593 18475 22627
rect 18417 22587 18475 22593
rect 18432 22556 18460 22587
rect 18598 22584 18604 22636
rect 18656 22624 18662 22636
rect 19260 22633 19288 22732
rect 19426 22720 19432 22732
rect 19484 22720 19490 22772
rect 22646 22760 22652 22772
rect 22607 22732 22652 22760
rect 22646 22720 22652 22732
rect 22704 22760 22710 22772
rect 23106 22760 23112 22772
rect 22704 22732 23112 22760
rect 22704 22720 22710 22732
rect 23106 22720 23112 22732
rect 23164 22720 23170 22772
rect 23198 22720 23204 22772
rect 23256 22760 23262 22772
rect 23750 22760 23756 22772
rect 23256 22732 23756 22760
rect 23256 22720 23262 22732
rect 23750 22720 23756 22732
rect 23808 22720 23814 22772
rect 25038 22720 25044 22772
rect 25096 22760 25102 22772
rect 25096 22732 25821 22760
rect 25096 22720 25102 22732
rect 24118 22692 24124 22704
rect 23492 22664 24124 22692
rect 23492 22636 23520 22664
rect 24118 22652 24124 22664
rect 24176 22652 24182 22704
rect 19061 22627 19119 22633
rect 19061 22624 19073 22627
rect 18656 22596 19073 22624
rect 18656 22584 18662 22596
rect 19061 22593 19073 22596
rect 19107 22593 19119 22627
rect 19061 22587 19119 22593
rect 19245 22627 19303 22633
rect 19245 22593 19257 22627
rect 19291 22593 19303 22627
rect 20254 22624 20260 22636
rect 20215 22596 20260 22624
rect 19245 22587 19303 22593
rect 20254 22584 20260 22596
rect 20312 22584 20318 22636
rect 20533 22627 20591 22633
rect 20533 22593 20545 22627
rect 20579 22624 20591 22627
rect 20714 22624 20720 22636
rect 20579 22596 20720 22624
rect 20579 22593 20591 22596
rect 20533 22587 20591 22593
rect 20714 22584 20720 22596
rect 20772 22584 20778 22636
rect 22738 22624 22744 22636
rect 22699 22596 22744 22624
rect 22738 22584 22744 22596
rect 22796 22584 22802 22636
rect 23474 22624 23480 22636
rect 23387 22596 23480 22624
rect 23474 22584 23480 22596
rect 23532 22584 23538 22636
rect 24489 22627 24547 22633
rect 24489 22624 24501 22627
rect 23860 22596 24501 22624
rect 23566 22556 23572 22568
rect 17092 22528 17137 22556
rect 17696 22528 18460 22556
rect 21284 22528 23428 22556
rect 23527 22528 23572 22556
rect 17092 22516 17098 22528
rect 18046 22488 18052 22500
rect 15344 22460 16528 22488
rect 16960 22460 18052 22488
rect 15344 22448 15350 22460
rect 16500 22432 16528 22460
rect 18046 22448 18052 22460
rect 18104 22448 18110 22500
rect 21284 22497 21312 22528
rect 21269 22491 21327 22497
rect 21269 22457 21281 22491
rect 21315 22457 21327 22491
rect 21269 22451 21327 22457
rect 22186 22448 22192 22500
rect 22244 22488 22250 22500
rect 22373 22491 22431 22497
rect 22373 22488 22385 22491
rect 22244 22460 22385 22488
rect 22244 22448 22250 22460
rect 22373 22457 22385 22460
rect 22419 22457 22431 22491
rect 23400 22488 23428 22528
rect 23566 22516 23572 22528
rect 23624 22516 23630 22568
rect 23860 22565 23888 22596
rect 24489 22593 24501 22596
rect 24535 22593 24547 22627
rect 24489 22587 24547 22593
rect 24578 22584 24584 22636
rect 24636 22624 24642 22636
rect 24762 22624 24768 22636
rect 24636 22596 24681 22624
rect 24723 22596 24768 22624
rect 24636 22584 24642 22596
rect 24762 22584 24768 22596
rect 24820 22584 24826 22636
rect 24857 22627 24915 22633
rect 24857 22593 24869 22627
rect 24903 22624 24915 22627
rect 25222 22624 25228 22636
rect 24903 22596 25228 22624
rect 24903 22593 24915 22596
rect 24857 22587 24915 22593
rect 25222 22584 25228 22596
rect 25280 22584 25286 22636
rect 25793 22633 25821 22732
rect 25866 22720 25872 22772
rect 25924 22760 25930 22772
rect 31018 22760 31024 22772
rect 25924 22732 31024 22760
rect 25924 22720 25930 22732
rect 31018 22720 31024 22732
rect 31076 22720 31082 22772
rect 33134 22760 33140 22772
rect 32140 22732 33140 22760
rect 27338 22692 27344 22704
rect 27299 22664 27344 22692
rect 27338 22652 27344 22664
rect 27396 22652 27402 22704
rect 28718 22652 28724 22704
rect 28776 22692 28782 22704
rect 31938 22692 31944 22704
rect 28776 22664 29868 22692
rect 28776 22652 28782 22664
rect 25685 22627 25743 22633
rect 25685 22593 25697 22627
rect 25731 22593 25743 22627
rect 25685 22587 25743 22593
rect 25777 22627 25835 22633
rect 25777 22593 25789 22627
rect 25823 22624 25835 22627
rect 26970 22624 26976 22636
rect 25823 22596 26976 22624
rect 25823 22593 25835 22596
rect 25777 22587 25835 22593
rect 23845 22559 23903 22565
rect 23845 22525 23857 22559
rect 23891 22525 23903 22559
rect 23845 22519 23903 22525
rect 24302 22516 24308 22568
rect 24360 22556 24366 22568
rect 25700 22556 25728 22587
rect 26970 22584 26976 22596
rect 27028 22584 27034 22636
rect 27062 22584 27068 22636
rect 27120 22624 27126 22636
rect 27522 22633 27528 22636
rect 27249 22627 27307 22633
rect 27120 22596 27165 22624
rect 27120 22584 27126 22596
rect 27249 22593 27261 22627
rect 27295 22593 27307 22627
rect 27249 22587 27307 22593
rect 27479 22627 27528 22633
rect 27479 22593 27491 22627
rect 27525 22593 27528 22627
rect 27479 22587 27528 22593
rect 26878 22556 26884 22568
rect 24360 22528 26884 22556
rect 24360 22516 24366 22528
rect 26878 22516 26884 22528
rect 26936 22516 26942 22568
rect 27264 22556 27292 22587
rect 27522 22584 27528 22587
rect 27580 22584 27586 22636
rect 28353 22627 28411 22633
rect 28353 22593 28365 22627
rect 28399 22593 28411 22627
rect 28534 22624 28540 22636
rect 28495 22596 28540 22624
rect 28353 22587 28411 22593
rect 27338 22556 27344 22568
rect 27264 22528 27344 22556
rect 27338 22516 27344 22528
rect 27396 22516 27402 22568
rect 28368 22556 28396 22587
rect 28534 22584 28540 22596
rect 28592 22584 28598 22636
rect 29086 22584 29092 22636
rect 29144 22624 29150 22636
rect 29181 22627 29239 22633
rect 29181 22624 29193 22627
rect 29144 22596 29193 22624
rect 29144 22584 29150 22596
rect 29181 22593 29193 22596
rect 29227 22593 29239 22627
rect 29362 22624 29368 22636
rect 29323 22596 29368 22624
rect 29181 22587 29239 22593
rect 28994 22556 29000 22568
rect 28368 22528 29000 22556
rect 28994 22516 29000 22528
rect 29052 22516 29058 22568
rect 29196 22556 29224 22587
rect 29362 22584 29368 22596
rect 29420 22584 29426 22636
rect 29840 22633 29868 22664
rect 31220 22664 31944 22692
rect 29825 22627 29883 22633
rect 29825 22593 29837 22627
rect 29871 22593 29883 22627
rect 29825 22587 29883 22593
rect 30009 22627 30067 22633
rect 30009 22593 30021 22627
rect 30055 22593 30067 22627
rect 30009 22587 30067 22593
rect 30024 22556 30052 22587
rect 30466 22584 30472 22636
rect 30524 22624 30530 22636
rect 31220 22633 31248 22664
rect 31938 22652 31944 22664
rect 31996 22652 32002 22704
rect 30561 22627 30619 22633
rect 30561 22624 30573 22627
rect 30524 22596 30573 22624
rect 30524 22584 30530 22596
rect 30561 22593 30573 22596
rect 30607 22593 30619 22627
rect 30561 22587 30619 22593
rect 30745 22627 30803 22633
rect 30745 22593 30757 22627
rect 30791 22593 30803 22627
rect 30745 22587 30803 22593
rect 31205 22627 31263 22633
rect 31205 22593 31217 22627
rect 31251 22593 31263 22627
rect 31205 22587 31263 22593
rect 31297 22627 31355 22633
rect 31297 22593 31309 22627
rect 31343 22624 31355 22627
rect 31386 22624 31392 22636
rect 31343 22596 31392 22624
rect 31343 22593 31355 22596
rect 31297 22587 31355 22593
rect 30650 22556 30656 22568
rect 29196 22528 30052 22556
rect 30484 22528 30656 22556
rect 30484 22488 30512 22528
rect 30650 22516 30656 22528
rect 30708 22516 30714 22568
rect 30760 22556 30788 22587
rect 31312 22556 31340 22587
rect 31386 22584 31392 22596
rect 31444 22584 31450 22636
rect 32140 22633 32168 22732
rect 33134 22720 33140 22732
rect 33192 22720 33198 22772
rect 34609 22763 34667 22769
rect 34609 22760 34621 22763
rect 33612 22732 34621 22760
rect 33612 22704 33640 22732
rect 34609 22729 34621 22732
rect 34655 22729 34667 22763
rect 34609 22723 34667 22729
rect 32217 22695 32275 22701
rect 32217 22661 32229 22695
rect 32263 22692 32275 22695
rect 33594 22692 33600 22704
rect 32263 22664 32996 22692
rect 33555 22664 33600 22692
rect 32263 22661 32275 22664
rect 32217 22655 32275 22661
rect 32125 22627 32183 22633
rect 32125 22593 32137 22627
rect 32171 22593 32183 22627
rect 32125 22587 32183 22593
rect 32309 22627 32367 22633
rect 32309 22593 32321 22627
rect 32355 22624 32367 22627
rect 32858 22624 32864 22636
rect 32355 22596 32864 22624
rect 32355 22593 32367 22596
rect 32309 22587 32367 22593
rect 32858 22584 32864 22596
rect 32916 22584 32922 22636
rect 32968 22633 32996 22664
rect 33594 22652 33600 22664
rect 33652 22652 33658 22704
rect 33813 22695 33871 22701
rect 33813 22661 33825 22695
rect 33859 22692 33871 22695
rect 34425 22695 34483 22701
rect 34425 22692 34437 22695
rect 33859 22664 34437 22692
rect 33859 22661 33871 22664
rect 33813 22655 33871 22661
rect 34425 22661 34437 22664
rect 34471 22692 34483 22695
rect 35618 22692 35624 22704
rect 34471 22664 35624 22692
rect 34471 22661 34483 22664
rect 34425 22655 34483 22661
rect 35618 22652 35624 22664
rect 35676 22652 35682 22704
rect 32953 22627 33011 22633
rect 32953 22593 32965 22627
rect 32999 22593 33011 22627
rect 32953 22587 33011 22593
rect 34701 22627 34759 22633
rect 34701 22593 34713 22627
rect 34747 22593 34759 22627
rect 34701 22587 34759 22593
rect 35345 22627 35403 22633
rect 35345 22593 35357 22627
rect 35391 22593 35403 22627
rect 35345 22587 35403 22593
rect 35437 22627 35495 22633
rect 35437 22593 35449 22627
rect 35483 22624 35495 22627
rect 36078 22624 36084 22636
rect 35483 22596 36084 22624
rect 35483 22593 35495 22596
rect 35437 22587 35495 22593
rect 31478 22556 31484 22568
rect 30760 22528 31340 22556
rect 31439 22528 31484 22556
rect 31478 22516 31484 22528
rect 31536 22516 31542 22568
rect 32769 22559 32827 22565
rect 32769 22525 32781 22559
rect 32815 22556 32827 22559
rect 33226 22556 33232 22568
rect 32815 22528 33232 22556
rect 32815 22525 32827 22528
rect 32769 22519 32827 22525
rect 33226 22516 33232 22528
rect 33284 22556 33290 22568
rect 33284 22528 33824 22556
rect 33284 22516 33290 22528
rect 23400 22460 30512 22488
rect 30561 22491 30619 22497
rect 22373 22451 22431 22457
rect 30561 22457 30573 22491
rect 30607 22488 30619 22491
rect 32122 22488 32128 22500
rect 30607 22460 32128 22488
rect 30607 22457 30619 22460
rect 30561 22451 30619 22457
rect 32122 22448 32128 22460
rect 32180 22448 32186 22500
rect 33594 22488 33600 22500
rect 33060 22460 33600 22488
rect 12124 22392 13124 22420
rect 12124 22380 12130 22392
rect 15378 22380 15384 22432
rect 15436 22420 15442 22432
rect 15565 22423 15623 22429
rect 15565 22420 15577 22423
rect 15436 22392 15577 22420
rect 15436 22380 15442 22392
rect 15565 22389 15577 22392
rect 15611 22389 15623 22423
rect 15565 22383 15623 22389
rect 16482 22380 16488 22432
rect 16540 22420 16546 22432
rect 18233 22423 18291 22429
rect 18233 22420 18245 22423
rect 16540 22392 18245 22420
rect 16540 22380 16546 22392
rect 18233 22389 18245 22392
rect 18279 22389 18291 22423
rect 18233 22383 18291 22389
rect 19429 22423 19487 22429
rect 19429 22389 19441 22423
rect 19475 22420 19487 22423
rect 20254 22420 20260 22432
rect 19475 22392 20260 22420
rect 19475 22389 19487 22392
rect 19429 22383 19487 22389
rect 20254 22380 20260 22392
rect 20312 22380 20318 22432
rect 22002 22420 22008 22432
rect 21963 22392 22008 22420
rect 22002 22380 22008 22392
rect 22060 22380 22066 22432
rect 22094 22380 22100 22432
rect 22152 22420 22158 22432
rect 22281 22423 22339 22429
rect 22281 22420 22293 22423
rect 22152 22392 22293 22420
rect 22152 22380 22158 22392
rect 22281 22389 22293 22392
rect 22327 22389 22339 22423
rect 22281 22383 22339 22389
rect 22465 22423 22523 22429
rect 22465 22389 22477 22423
rect 22511 22420 22523 22423
rect 22646 22420 22652 22432
rect 22511 22392 22652 22420
rect 22511 22389 22523 22392
rect 22465 22383 22523 22389
rect 22646 22380 22652 22392
rect 22704 22380 22710 22432
rect 24305 22423 24363 22429
rect 24305 22389 24317 22423
rect 24351 22420 24363 22423
rect 25866 22420 25872 22432
rect 24351 22392 25872 22420
rect 24351 22389 24363 22392
rect 24305 22383 24363 22389
rect 25866 22380 25872 22392
rect 25924 22380 25930 22432
rect 26786 22380 26792 22432
rect 26844 22420 26850 22432
rect 27522 22420 27528 22432
rect 26844 22392 27528 22420
rect 26844 22380 26850 22392
rect 27522 22380 27528 22392
rect 27580 22380 27586 22432
rect 27617 22423 27675 22429
rect 27617 22389 27629 22423
rect 27663 22420 27675 22423
rect 27798 22420 27804 22432
rect 27663 22392 27804 22420
rect 27663 22389 27675 22392
rect 27617 22383 27675 22389
rect 27798 22380 27804 22392
rect 27856 22380 27862 22432
rect 28258 22380 28264 22432
rect 28316 22420 28322 22432
rect 28718 22420 28724 22432
rect 28316 22392 28724 22420
rect 28316 22380 28322 22392
rect 28718 22380 28724 22392
rect 28776 22380 28782 22432
rect 28994 22380 29000 22432
rect 29052 22420 29058 22432
rect 29273 22423 29331 22429
rect 29273 22420 29285 22423
rect 29052 22392 29285 22420
rect 29052 22380 29058 22392
rect 29273 22389 29285 22392
rect 29319 22389 29331 22423
rect 29914 22420 29920 22432
rect 29875 22392 29920 22420
rect 29273 22383 29331 22389
rect 29914 22380 29920 22392
rect 29972 22380 29978 22432
rect 31389 22423 31447 22429
rect 31389 22389 31401 22423
rect 31435 22420 31447 22423
rect 33060 22420 33088 22460
rect 33594 22448 33600 22460
rect 33652 22448 33658 22500
rect 33796 22488 33824 22528
rect 34716 22488 34744 22587
rect 33796 22460 34744 22488
rect 35360 22488 35388 22587
rect 36078 22584 36084 22596
rect 36136 22584 36142 22636
rect 36262 22624 36268 22636
rect 36223 22596 36268 22624
rect 36262 22584 36268 22596
rect 36320 22584 36326 22636
rect 35621 22559 35679 22565
rect 35621 22525 35633 22559
rect 35667 22556 35679 22559
rect 36280 22556 36308 22584
rect 35667 22528 36308 22556
rect 35667 22525 35679 22528
rect 35621 22519 35679 22525
rect 35360 22460 35756 22488
rect 31435 22392 33088 22420
rect 33137 22423 33195 22429
rect 31435 22389 31447 22392
rect 31389 22383 31447 22389
rect 33137 22389 33149 22423
rect 33183 22420 33195 22423
rect 33226 22420 33232 22432
rect 33183 22392 33232 22420
rect 33183 22389 33195 22392
rect 33137 22383 33195 22389
rect 33226 22380 33232 22392
rect 33284 22380 33290 22432
rect 33796 22429 33824 22460
rect 33781 22423 33839 22429
rect 33781 22389 33793 22423
rect 33827 22389 33839 22423
rect 33962 22420 33968 22432
rect 33923 22392 33968 22420
rect 33781 22383 33839 22389
rect 33962 22380 33968 22392
rect 34020 22380 34026 22432
rect 34422 22420 34428 22432
rect 34383 22392 34428 22420
rect 34422 22380 34428 22392
rect 34480 22380 34486 22432
rect 35526 22380 35532 22432
rect 35584 22420 35590 22432
rect 35728 22420 35756 22460
rect 35894 22448 35900 22500
rect 35952 22488 35958 22500
rect 36449 22491 36507 22497
rect 36449 22488 36461 22491
rect 35952 22460 36461 22488
rect 35952 22448 35958 22460
rect 36449 22457 36461 22460
rect 36495 22488 36507 22491
rect 36630 22488 36636 22500
rect 36495 22460 36636 22488
rect 36495 22457 36507 22460
rect 36449 22451 36507 22457
rect 36630 22448 36636 22460
rect 36688 22448 36694 22500
rect 36265 22423 36323 22429
rect 36265 22420 36277 22423
rect 35584 22392 35629 22420
rect 35728 22392 36277 22420
rect 35584 22380 35590 22392
rect 36265 22389 36277 22392
rect 36311 22420 36323 22423
rect 36722 22420 36728 22432
rect 36311 22392 36728 22420
rect 36311 22389 36323 22392
rect 36265 22383 36323 22389
rect 36722 22380 36728 22392
rect 36780 22380 36786 22432
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 14458 22176 14464 22228
rect 14516 22216 14522 22228
rect 14829 22219 14887 22225
rect 14829 22216 14841 22219
rect 14516 22188 14841 22216
rect 14516 22176 14522 22188
rect 14829 22185 14841 22188
rect 14875 22185 14887 22219
rect 17770 22216 17776 22228
rect 14829 22179 14887 22185
rect 15580 22188 17776 22216
rect 11146 22148 11152 22160
rect 11107 22120 11152 22148
rect 11146 22108 11152 22120
rect 11204 22108 11210 22160
rect 15194 22108 15200 22160
rect 15252 22148 15258 22160
rect 15470 22148 15476 22160
rect 15252 22120 15476 22148
rect 15252 22108 15258 22120
rect 15470 22108 15476 22120
rect 15528 22108 15534 22160
rect 9493 22083 9551 22089
rect 9493 22049 9505 22083
rect 9539 22080 9551 22083
rect 9674 22080 9680 22092
rect 9539 22052 9680 22080
rect 9539 22049 9551 22052
rect 9493 22043 9551 22049
rect 9674 22040 9680 22052
rect 9732 22040 9738 22092
rect 9950 22080 9956 22092
rect 9911 22052 9956 22080
rect 9950 22040 9956 22052
rect 10008 22040 10014 22092
rect 13078 22080 13084 22092
rect 12176 22052 13084 22080
rect 1394 22012 1400 22024
rect 1355 21984 1400 22012
rect 1394 21972 1400 21984
rect 1452 21972 1458 22024
rect 8846 21972 8852 22024
rect 8904 22012 8910 22024
rect 9585 22015 9643 22021
rect 9585 22012 9597 22015
rect 8904 21984 9597 22012
rect 8904 21972 8910 21984
rect 9585 21981 9597 21984
rect 9631 21981 9643 22015
rect 9585 21975 9643 21981
rect 11606 21972 11612 22024
rect 11664 22012 11670 22024
rect 11971 22021 11977 22024
rect 11865 22015 11923 22021
rect 11865 22012 11877 22015
rect 11664 21984 11877 22012
rect 11664 21972 11670 21984
rect 10962 21944 10968 21956
rect 10923 21916 10968 21944
rect 10962 21904 10968 21916
rect 11020 21904 11026 21956
rect 1581 21879 1639 21885
rect 1581 21845 1593 21879
rect 1627 21876 1639 21879
rect 7926 21876 7932 21888
rect 1627 21848 7932 21876
rect 1627 21845 1639 21848
rect 1581 21839 1639 21845
rect 7926 21836 7932 21848
rect 7984 21836 7990 21888
rect 11609 21879 11667 21885
rect 11609 21845 11621 21879
rect 11655 21876 11667 21879
rect 11698 21876 11704 21888
rect 11655 21848 11704 21876
rect 11655 21845 11667 21848
rect 11609 21839 11667 21845
rect 11698 21836 11704 21848
rect 11756 21836 11762 21888
rect 11808 21876 11836 21984
rect 11865 21981 11877 21984
rect 11911 21981 11923 22015
rect 11865 21975 11923 21981
rect 11958 22015 11977 22021
rect 11958 21981 11970 22015
rect 11958 21975 11977 21981
rect 11971 21972 11977 21975
rect 12029 21972 12035 22024
rect 12090 22015 12148 22021
rect 12090 21981 12102 22015
rect 12136 22012 12148 22015
rect 12176 22012 12204 22052
rect 13078 22040 13084 22052
rect 13136 22040 13142 22092
rect 15580 22080 15608 22188
rect 17770 22176 17776 22188
rect 17828 22176 17834 22228
rect 20714 22216 20720 22228
rect 20675 22188 20720 22216
rect 20714 22176 20720 22188
rect 20772 22176 20778 22228
rect 21637 22219 21695 22225
rect 21637 22185 21649 22219
rect 21683 22185 21695 22219
rect 22646 22216 22652 22228
rect 22607 22188 22652 22216
rect 21637 22179 21695 22185
rect 15654 22108 15660 22160
rect 15712 22148 15718 22160
rect 21652 22148 21680 22179
rect 22646 22176 22652 22188
rect 22704 22176 22710 22228
rect 22738 22176 22744 22228
rect 22796 22216 22802 22228
rect 23017 22219 23075 22225
rect 23017 22216 23029 22219
rect 22796 22188 23029 22216
rect 22796 22176 22802 22188
rect 23017 22185 23029 22188
rect 23063 22185 23075 22219
rect 23658 22216 23664 22228
rect 23619 22188 23664 22216
rect 23017 22179 23075 22185
rect 23658 22176 23664 22188
rect 23716 22176 23722 22228
rect 25314 22176 25320 22228
rect 25372 22216 25378 22228
rect 26050 22216 26056 22228
rect 25372 22188 26056 22216
rect 25372 22176 25378 22188
rect 26050 22176 26056 22188
rect 26108 22176 26114 22228
rect 26234 22216 26240 22228
rect 26195 22188 26240 22216
rect 26234 22176 26240 22188
rect 26292 22176 26298 22228
rect 28166 22176 28172 22228
rect 28224 22216 28230 22228
rect 28442 22216 28448 22228
rect 28224 22188 28448 22216
rect 28224 22176 28230 22188
rect 28442 22176 28448 22188
rect 28500 22216 28506 22228
rect 30558 22216 30564 22228
rect 28500 22188 30420 22216
rect 30519 22188 30564 22216
rect 28500 22176 28506 22188
rect 24394 22148 24400 22160
rect 15712 22120 19012 22148
rect 21652 22120 24400 22148
rect 15712 22108 15718 22120
rect 16390 22080 16396 22092
rect 14200 22052 15608 22080
rect 16351 22052 16396 22080
rect 12136 21984 12204 22012
rect 12136 21981 12148 21984
rect 12090 21975 12148 21981
rect 12250 21972 12256 22024
rect 12308 22012 12314 22024
rect 13541 22015 13599 22021
rect 12308 21984 12353 22012
rect 12308 21972 12314 21984
rect 13541 21981 13553 22015
rect 13587 22012 13599 22015
rect 14090 22012 14096 22024
rect 13587 21984 14096 22012
rect 13587 21981 13599 21984
rect 13541 21975 13599 21981
rect 14090 21972 14096 21984
rect 14148 21972 14154 22024
rect 14200 22021 14228 22052
rect 16390 22040 16396 22052
rect 16448 22080 16454 22092
rect 16448 22052 17468 22080
rect 16448 22040 16454 22052
rect 14185 22015 14243 22021
rect 14185 21981 14197 22015
rect 14231 21981 14243 22015
rect 14185 21975 14243 21981
rect 14369 22015 14427 22021
rect 14369 21981 14381 22015
rect 14415 21981 14427 22015
rect 14369 21975 14427 21981
rect 15013 22015 15071 22021
rect 15013 21981 15025 22015
rect 15059 22012 15071 22015
rect 15194 22012 15200 22024
rect 15059 21984 15200 22012
rect 15059 21981 15071 21984
rect 15013 21975 15071 21981
rect 14384 21944 14412 21975
rect 15194 21972 15200 21984
rect 15252 21972 15258 22024
rect 15473 22015 15531 22021
rect 15473 21981 15485 22015
rect 15519 21981 15531 22015
rect 15654 22012 15660 22024
rect 15615 21984 15660 22012
rect 15473 21975 15531 21981
rect 15378 21944 15384 21956
rect 14384 21916 15384 21944
rect 15378 21904 15384 21916
rect 15436 21904 15442 21956
rect 15488 21944 15516 21975
rect 15654 21972 15660 21984
rect 15712 21972 15718 22024
rect 15930 21972 15936 22024
rect 15988 22012 15994 22024
rect 17440 22021 17468 22052
rect 16117 22015 16175 22021
rect 16117 22012 16129 22015
rect 15988 21984 16129 22012
rect 15988 21972 15994 21984
rect 16117 21981 16129 21984
rect 16163 21981 16175 22015
rect 16117 21975 16175 21981
rect 17405 22015 17468 22021
rect 17405 21981 17417 22015
rect 17451 21986 17468 22015
rect 17770 22012 17776 22024
rect 17451 21981 17463 21986
rect 17731 21984 17776 22012
rect 17405 21975 17463 21981
rect 17770 21972 17776 21984
rect 17828 21972 17834 22024
rect 18230 21972 18236 22024
rect 18288 22012 18294 22024
rect 18693 22015 18751 22021
rect 18693 22012 18705 22015
rect 18288 21984 18705 22012
rect 18288 21972 18294 21984
rect 18693 21981 18705 21984
rect 18739 21981 18751 22015
rect 18984 22012 19012 22120
rect 24394 22108 24400 22120
rect 24452 22108 24458 22160
rect 24670 22108 24676 22160
rect 24728 22148 24734 22160
rect 24728 22120 25084 22148
rect 24728 22108 24734 22120
rect 20346 22040 20352 22092
rect 20404 22080 20410 22092
rect 23106 22080 23112 22092
rect 20404 22052 22094 22080
rect 23067 22052 23112 22080
rect 20404 22040 20410 22052
rect 19058 22012 19064 22024
rect 18984 21984 19064 22012
rect 18693 21975 18751 21981
rect 19058 21972 19064 21984
rect 19116 22012 19122 22024
rect 19245 22015 19303 22021
rect 19245 22012 19257 22015
rect 19116 21984 19257 22012
rect 19116 21972 19122 21984
rect 19245 21981 19257 21984
rect 19291 21981 19303 22015
rect 19426 22012 19432 22024
rect 19387 21984 19432 22012
rect 19245 21975 19303 21981
rect 19426 21972 19432 21984
rect 19484 21972 19490 22024
rect 20254 22012 20260 22024
rect 20215 21984 20260 22012
rect 20254 21972 20260 21984
rect 20312 21972 20318 22024
rect 20901 22015 20959 22021
rect 20901 21981 20913 22015
rect 20947 21981 20959 22015
rect 22066 22012 22094 22052
rect 23106 22040 23112 22052
rect 23164 22040 23170 22092
rect 23658 22080 23664 22092
rect 23400 22052 23664 22080
rect 22833 22015 22891 22021
rect 22066 21984 22784 22012
rect 20901 21975 20959 21981
rect 16942 21944 16948 21956
rect 15488 21916 16948 21944
rect 16942 21904 16948 21916
rect 17000 21904 17006 21956
rect 17589 21947 17647 21953
rect 17589 21944 17601 21947
rect 17052 21916 17601 21944
rect 13078 21876 13084 21888
rect 11808 21848 13084 21876
rect 13078 21836 13084 21848
rect 13136 21836 13142 21888
rect 13354 21876 13360 21888
rect 13315 21848 13360 21876
rect 13354 21836 13360 21848
rect 13412 21836 13418 21888
rect 14369 21879 14427 21885
rect 14369 21845 14381 21879
rect 14415 21876 14427 21879
rect 16298 21876 16304 21888
rect 14415 21848 16304 21876
rect 14415 21845 14427 21848
rect 14369 21839 14427 21845
rect 16298 21836 16304 21848
rect 16356 21876 16362 21888
rect 17052 21876 17080 21916
rect 17589 21913 17601 21916
rect 17635 21913 17647 21947
rect 17589 21907 17647 21913
rect 17678 21904 17684 21956
rect 17736 21944 17742 21956
rect 19613 21947 19671 21953
rect 17736 21916 17781 21944
rect 17736 21904 17742 21916
rect 19613 21913 19625 21947
rect 19659 21944 19671 21947
rect 20916 21944 20944 21975
rect 19659 21916 20944 21944
rect 21453 21947 21511 21953
rect 19659 21913 19671 21916
rect 19613 21907 19671 21913
rect 21453 21913 21465 21947
rect 21499 21944 21511 21947
rect 21542 21944 21548 21956
rect 21499 21916 21548 21944
rect 21499 21913 21511 21916
rect 21453 21907 21511 21913
rect 21542 21904 21548 21916
rect 21600 21904 21606 21956
rect 21669 21947 21727 21953
rect 21669 21913 21681 21947
rect 21715 21944 21727 21947
rect 22002 21944 22008 21956
rect 21715 21916 22008 21944
rect 21715 21913 21727 21916
rect 21669 21907 21727 21913
rect 22002 21904 22008 21916
rect 22060 21904 22066 21956
rect 22756 21944 22784 21984
rect 22833 21981 22845 22015
rect 22879 22012 22891 22015
rect 23400 22012 23428 22052
rect 23658 22040 23664 22052
rect 23716 22040 23722 22092
rect 23842 22080 23848 22092
rect 23803 22052 23848 22080
rect 23842 22040 23848 22052
rect 23900 22080 23906 22092
rect 24946 22080 24952 22092
rect 23900 22052 24440 22080
rect 24907 22052 24952 22080
rect 23900 22040 23906 22052
rect 22879 21984 23428 22012
rect 22879 21981 22891 21984
rect 22833 21975 22891 21981
rect 23474 21972 23480 22024
rect 23532 22012 23538 22024
rect 24412 22021 24440 22052
rect 24946 22040 24952 22052
rect 25004 22040 25010 22092
rect 25056 22080 25084 22120
rect 26510 22108 26516 22160
rect 26568 22148 26574 22160
rect 26878 22148 26884 22160
rect 26568 22120 26884 22148
rect 26568 22108 26574 22120
rect 26878 22108 26884 22120
rect 26936 22108 26942 22160
rect 26973 22151 27031 22157
rect 26973 22117 26985 22151
rect 27019 22148 27031 22151
rect 27706 22148 27712 22160
rect 27019 22120 27712 22148
rect 27019 22117 27031 22120
rect 26973 22111 27031 22117
rect 27706 22108 27712 22120
rect 27764 22108 27770 22160
rect 28534 22108 28540 22160
rect 28592 22148 28598 22160
rect 29822 22148 29828 22160
rect 28592 22120 29828 22148
rect 28592 22108 28598 22120
rect 29822 22108 29828 22120
rect 29880 22108 29886 22160
rect 30392 22148 30420 22188
rect 30558 22176 30564 22188
rect 30616 22176 30622 22228
rect 33137 22219 33195 22225
rect 33137 22185 33149 22219
rect 33183 22216 33195 22219
rect 34606 22216 34612 22228
rect 33183 22188 34612 22216
rect 33183 22185 33195 22188
rect 33137 22179 33195 22185
rect 34606 22176 34612 22188
rect 34664 22176 34670 22228
rect 35529 22219 35587 22225
rect 35529 22185 35541 22219
rect 35575 22216 35587 22219
rect 35618 22216 35624 22228
rect 35575 22188 35624 22216
rect 35575 22185 35587 22188
rect 35529 22179 35587 22185
rect 35618 22176 35624 22188
rect 35676 22176 35682 22228
rect 33410 22148 33416 22160
rect 30392 22120 33416 22148
rect 33410 22108 33416 22120
rect 33468 22108 33474 22160
rect 33505 22151 33563 22157
rect 33505 22117 33517 22151
rect 33551 22148 33563 22151
rect 33686 22148 33692 22160
rect 33551 22120 33692 22148
rect 33551 22117 33563 22120
rect 33505 22111 33563 22117
rect 33686 22108 33692 22120
rect 33744 22108 33750 22160
rect 33778 22108 33784 22160
rect 33836 22148 33842 22160
rect 34793 22151 34851 22157
rect 34793 22148 34805 22151
rect 33836 22120 34805 22148
rect 33836 22108 33842 22120
rect 34793 22117 34805 22120
rect 34839 22117 34851 22151
rect 34793 22111 34851 22117
rect 25133 22083 25191 22089
rect 25133 22080 25145 22083
rect 25056 22052 25145 22080
rect 25133 22049 25145 22052
rect 25179 22049 25191 22083
rect 25133 22043 25191 22049
rect 26160 22052 27016 22080
rect 23569 22015 23627 22021
rect 23569 22012 23581 22015
rect 23532 21984 23581 22012
rect 23532 21972 23538 21984
rect 23569 21981 23581 21984
rect 23615 21981 23627 22015
rect 23569 21975 23627 21981
rect 24397 22015 24455 22021
rect 24397 21981 24409 22015
rect 24443 21981 24455 22015
rect 24397 21975 24455 21981
rect 24578 21972 24584 22024
rect 24636 22012 24642 22024
rect 24854 22012 24860 22024
rect 24636 21984 24860 22012
rect 24636 21972 24642 21984
rect 24854 21972 24860 21984
rect 24912 21972 24918 22024
rect 25225 22015 25283 22021
rect 25225 21981 25237 22015
rect 25271 21981 25283 22015
rect 25225 21975 25283 21981
rect 25240 21944 25268 21975
rect 25406 21972 25412 22024
rect 25464 22012 25470 22024
rect 26160 22021 26188 22052
rect 26145 22015 26203 22021
rect 26145 22012 26157 22015
rect 25464 21984 26157 22012
rect 25464 21972 25470 21984
rect 26145 21981 26157 21984
rect 26191 21981 26203 22015
rect 26145 21975 26203 21981
rect 26881 22015 26939 22021
rect 26881 21981 26893 22015
rect 26927 21981 26939 22015
rect 26988 22012 27016 22052
rect 27062 22040 27068 22092
rect 27120 22080 27126 22092
rect 27157 22083 27215 22089
rect 27157 22080 27169 22083
rect 27120 22052 27169 22080
rect 27120 22040 27126 22052
rect 27157 22049 27169 22052
rect 27203 22049 27215 22083
rect 27157 22043 27215 22049
rect 27522 22040 27528 22092
rect 27580 22080 27586 22092
rect 28077 22083 28135 22089
rect 28077 22080 28089 22083
rect 27580 22052 28089 22080
rect 27580 22040 27586 22052
rect 28077 22049 28089 22052
rect 28123 22049 28135 22083
rect 28258 22080 28264 22092
rect 28219 22052 28264 22080
rect 28077 22043 28135 22049
rect 28258 22040 28264 22052
rect 28316 22040 28322 22092
rect 28353 22083 28411 22089
rect 28353 22049 28365 22083
rect 28399 22080 28411 22083
rect 28399 22052 30328 22080
rect 28399 22049 28411 22052
rect 28353 22043 28411 22049
rect 27982 22012 27988 22024
rect 26988 21984 27988 22012
rect 26881 21975 26939 21981
rect 22756 21916 25268 21944
rect 26896 21944 26924 21975
rect 27982 21972 27988 21984
rect 28040 21972 28046 22024
rect 28169 22015 28227 22021
rect 28169 21981 28181 22015
rect 28215 21981 28227 22015
rect 28169 21975 28227 21981
rect 28184 21944 28212 21975
rect 28994 21972 29000 22024
rect 29052 22012 29058 22024
rect 29546 22012 29552 22024
rect 29052 21984 29552 22012
rect 29052 21972 29058 21984
rect 29546 21972 29552 21984
rect 29604 21972 29610 22024
rect 29733 22015 29791 22021
rect 29733 21981 29745 22015
rect 29779 22012 29791 22015
rect 29822 22012 29828 22024
rect 29779 21984 29828 22012
rect 29779 21981 29791 21984
rect 29733 21975 29791 21981
rect 29822 21972 29828 21984
rect 29880 21972 29886 22024
rect 30193 22015 30251 22021
rect 30193 21981 30205 22015
rect 30239 21981 30251 22015
rect 30300 22012 30328 22052
rect 30742 22040 30748 22092
rect 30800 22080 30806 22092
rect 31570 22080 31576 22092
rect 30800 22052 31576 22080
rect 30800 22040 30806 22052
rect 31570 22040 31576 22052
rect 31628 22040 31634 22092
rect 32490 22040 32496 22092
rect 32548 22080 32554 22092
rect 33597 22083 33655 22089
rect 33597 22080 33609 22083
rect 32548 22052 33609 22080
rect 32548 22040 32554 22052
rect 33597 22049 33609 22052
rect 33643 22080 33655 22083
rect 34977 22083 35035 22089
rect 34977 22080 34989 22083
rect 33643 22052 34989 22080
rect 33643 22049 33655 22052
rect 33597 22043 33655 22049
rect 34977 22049 34989 22052
rect 35023 22049 35035 22083
rect 34977 22043 35035 22049
rect 31202 22012 31208 22024
rect 30300 21984 30788 22012
rect 31163 21984 31208 22012
rect 30193 21975 30251 21981
rect 29641 21947 29699 21953
rect 29641 21944 29653 21947
rect 26896 21916 28120 21944
rect 28184 21916 29653 21944
rect 16356 21848 17080 21876
rect 16356 21836 16362 21848
rect 17126 21836 17132 21888
rect 17184 21876 17190 21888
rect 17957 21879 18015 21885
rect 17957 21876 17969 21879
rect 17184 21848 17969 21876
rect 17184 21836 17190 21848
rect 17957 21845 17969 21848
rect 18003 21845 18015 21879
rect 17957 21839 18015 21845
rect 18138 21836 18144 21888
rect 18196 21876 18202 21888
rect 18509 21879 18567 21885
rect 18509 21876 18521 21879
rect 18196 21848 18521 21876
rect 18196 21836 18202 21848
rect 18509 21845 18521 21848
rect 18555 21845 18567 21879
rect 18509 21839 18567 21845
rect 20073 21879 20131 21885
rect 20073 21845 20085 21879
rect 20119 21876 20131 21879
rect 20806 21876 20812 21888
rect 20119 21848 20812 21876
rect 20119 21845 20131 21848
rect 20073 21839 20131 21845
rect 20806 21836 20812 21848
rect 20864 21836 20870 21888
rect 21818 21876 21824 21888
rect 21779 21848 21824 21876
rect 21818 21836 21824 21848
rect 21876 21836 21882 21888
rect 23474 21836 23480 21888
rect 23532 21876 23538 21888
rect 23845 21879 23903 21885
rect 23845 21876 23857 21879
rect 23532 21848 23857 21876
rect 23532 21836 23538 21848
rect 23845 21845 23857 21848
rect 23891 21845 23903 21879
rect 23845 21839 23903 21845
rect 24489 21879 24547 21885
rect 24489 21845 24501 21879
rect 24535 21876 24547 21879
rect 26142 21876 26148 21888
rect 24535 21848 26148 21876
rect 24535 21845 24547 21848
rect 24489 21839 24547 21845
rect 26142 21836 26148 21848
rect 26200 21836 26206 21888
rect 27154 21876 27160 21888
rect 27115 21848 27160 21876
rect 27154 21836 27160 21848
rect 27212 21836 27218 21888
rect 27890 21876 27896 21888
rect 27851 21848 27896 21876
rect 27890 21836 27896 21848
rect 27948 21836 27954 21888
rect 28092 21876 28120 21916
rect 29641 21913 29653 21916
rect 29687 21913 29699 21947
rect 30208 21944 30236 21975
rect 30650 21944 30656 21956
rect 30208 21916 30656 21944
rect 29641 21907 29699 21913
rect 30650 21904 30656 21916
rect 30708 21904 30714 21956
rect 28534 21876 28540 21888
rect 28092 21848 28540 21876
rect 28534 21836 28540 21848
rect 28592 21836 28598 21888
rect 28718 21836 28724 21888
rect 28776 21876 28782 21888
rect 30006 21876 30012 21888
rect 28776 21848 30012 21876
rect 28776 21836 28782 21848
rect 30006 21836 30012 21848
rect 30064 21836 30070 21888
rect 30098 21836 30104 21888
rect 30156 21876 30162 21888
rect 30760 21885 30788 21984
rect 31202 21972 31208 21984
rect 31260 21972 31266 22024
rect 31389 22015 31447 22021
rect 31389 21981 31401 22015
rect 31435 22012 31447 22015
rect 32214 22012 32220 22024
rect 31435 21984 32220 22012
rect 31435 21981 31447 21984
rect 31389 21975 31447 21981
rect 32214 21972 32220 21984
rect 32272 22012 32278 22024
rect 32401 22015 32459 22021
rect 32401 22012 32413 22015
rect 32272 21984 32413 22012
rect 32272 21972 32278 21984
rect 32401 21981 32413 21984
rect 32447 21981 32459 22015
rect 32401 21975 32459 21981
rect 33321 22015 33379 22021
rect 33321 21981 33333 22015
rect 33367 22012 33379 22015
rect 34054 22012 34060 22024
rect 33367 21984 34060 22012
rect 33367 21981 33379 21984
rect 33321 21975 33379 21981
rect 34054 21972 34060 21984
rect 34112 22012 34118 22024
rect 34701 22015 34759 22021
rect 34701 22012 34713 22015
rect 34112 21984 34713 22012
rect 34112 21972 34118 21984
rect 34701 21981 34713 21984
rect 34747 21981 34759 22015
rect 35434 22012 35440 22024
rect 35395 21984 35440 22012
rect 34701 21975 34759 21981
rect 35434 21972 35440 21984
rect 35492 21972 35498 22024
rect 35618 22012 35624 22024
rect 35579 21984 35624 22012
rect 35618 21972 35624 21984
rect 35676 21972 35682 22024
rect 37366 22012 37372 22024
rect 37327 21984 37372 22012
rect 37366 21972 37372 21984
rect 37424 21972 37430 22024
rect 37734 22012 37740 22024
rect 37695 21984 37740 22012
rect 37734 21972 37740 21984
rect 37792 21972 37798 22024
rect 30561 21879 30619 21885
rect 30561 21876 30573 21879
rect 30156 21848 30573 21876
rect 30156 21836 30162 21848
rect 30561 21845 30573 21848
rect 30607 21845 30619 21879
rect 30561 21839 30619 21845
rect 30745 21879 30803 21885
rect 30745 21845 30757 21879
rect 30791 21845 30803 21879
rect 30745 21839 30803 21845
rect 30834 21836 30840 21888
rect 30892 21876 30898 21888
rect 31297 21879 31355 21885
rect 31297 21876 31309 21879
rect 30892 21848 31309 21876
rect 30892 21836 30898 21848
rect 31297 21845 31309 21848
rect 31343 21845 31355 21879
rect 32490 21876 32496 21888
rect 32451 21848 32496 21876
rect 31297 21839 31355 21845
rect 32490 21836 32496 21848
rect 32548 21836 32554 21888
rect 34698 21876 34704 21888
rect 34659 21848 34704 21876
rect 34698 21836 34704 21848
rect 34756 21836 34762 21888
rect 38102 21876 38108 21888
rect 38063 21848 38108 21876
rect 38102 21836 38108 21848
rect 38160 21836 38166 21888
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 8665 21675 8723 21681
rect 8665 21641 8677 21675
rect 8711 21672 8723 21675
rect 8846 21672 8852 21684
rect 8711 21644 8852 21672
rect 8711 21641 8723 21644
rect 8665 21635 8723 21641
rect 8846 21632 8852 21644
rect 8904 21632 8910 21684
rect 10042 21632 10048 21684
rect 10100 21672 10106 21684
rect 10226 21672 10232 21684
rect 10100 21644 10232 21672
rect 10100 21632 10106 21644
rect 10226 21632 10232 21644
rect 10284 21672 10290 21684
rect 10597 21675 10655 21681
rect 10597 21672 10609 21675
rect 10284 21644 10609 21672
rect 10284 21632 10290 21644
rect 10597 21641 10609 21644
rect 10643 21641 10655 21675
rect 12618 21672 12624 21684
rect 10597 21635 10655 21641
rect 12406 21644 12624 21672
rect 7552 21539 7610 21545
rect 7552 21505 7564 21539
rect 7598 21536 7610 21539
rect 8864 21536 8892 21632
rect 9309 21607 9367 21613
rect 9309 21573 9321 21607
rect 9355 21604 9367 21607
rect 9766 21604 9772 21616
rect 9355 21576 9772 21604
rect 9355 21573 9367 21576
rect 9309 21567 9367 21573
rect 9766 21564 9772 21576
rect 9824 21564 9830 21616
rect 12406 21604 12434 21644
rect 12618 21632 12624 21644
rect 12676 21672 12682 21684
rect 13446 21672 13452 21684
rect 12676 21644 13452 21672
rect 12676 21632 12682 21644
rect 13446 21632 13452 21644
rect 13504 21632 13510 21684
rect 14366 21672 14372 21684
rect 14279 21644 14372 21672
rect 14366 21632 14372 21644
rect 14424 21672 14430 21684
rect 18141 21675 18199 21681
rect 14424 21644 17632 21672
rect 14424 21632 14430 21644
rect 13170 21604 13176 21616
rect 12268 21576 12434 21604
rect 13004 21576 13176 21604
rect 12268 21545 12296 21576
rect 9677 21539 9735 21545
rect 9677 21536 9689 21539
rect 7598 21508 8800 21536
rect 8864 21508 9689 21536
rect 7598 21505 7610 21508
rect 7552 21499 7610 21505
rect 7006 21428 7012 21480
rect 7064 21468 7070 21480
rect 7282 21468 7288 21480
rect 7064 21440 7288 21468
rect 7064 21428 7070 21440
rect 7282 21428 7288 21440
rect 7340 21428 7346 21480
rect 8772 21400 8800 21508
rect 9677 21505 9689 21508
rect 9723 21536 9735 21539
rect 10505 21539 10563 21545
rect 10505 21536 10517 21539
rect 9723 21508 10517 21536
rect 9723 21505 9735 21508
rect 9677 21499 9735 21505
rect 10505 21505 10517 21508
rect 10551 21505 10563 21539
rect 10505 21499 10563 21505
rect 12161 21539 12219 21545
rect 12161 21505 12173 21539
rect 12207 21505 12219 21539
rect 12161 21499 12219 21505
rect 12253 21539 12311 21545
rect 12253 21505 12265 21539
rect 12299 21505 12311 21539
rect 12253 21499 12311 21505
rect 12437 21539 12495 21545
rect 12437 21505 12449 21539
rect 12483 21536 12495 21539
rect 12618 21536 12624 21548
rect 12483 21508 12624 21536
rect 12483 21505 12495 21508
rect 12437 21499 12495 21505
rect 9769 21471 9827 21477
rect 9769 21437 9781 21471
rect 9815 21468 9827 21471
rect 11146 21468 11152 21480
rect 9815 21440 11152 21468
rect 9815 21437 9827 21440
rect 9769 21431 9827 21437
rect 11146 21428 11152 21440
rect 11204 21428 11210 21480
rect 12176 21468 12204 21499
rect 12618 21496 12624 21508
rect 12676 21496 12682 21548
rect 13004 21545 13032 21576
rect 13170 21564 13176 21576
rect 13228 21564 13234 21616
rect 15378 21604 15384 21616
rect 15339 21576 15384 21604
rect 15378 21564 15384 21576
rect 15436 21564 15442 21616
rect 13262 21545 13268 21548
rect 12989 21539 13047 21545
rect 12989 21505 13001 21539
rect 13035 21505 13047 21539
rect 12989 21499 13047 21505
rect 13256 21499 13268 21545
rect 13320 21536 13326 21548
rect 15289 21539 15347 21545
rect 13320 21508 13356 21536
rect 13262 21496 13268 21499
rect 13320 21496 13326 21508
rect 15289 21505 15301 21539
rect 15335 21536 15347 21539
rect 15470 21536 15476 21548
rect 15335 21508 15476 21536
rect 15335 21505 15347 21508
rect 15289 21499 15347 21505
rect 15470 21496 15476 21508
rect 15528 21496 15534 21548
rect 15930 21536 15936 21548
rect 15891 21508 15936 21536
rect 15930 21496 15936 21508
rect 15988 21496 15994 21548
rect 16114 21536 16120 21548
rect 16075 21508 16120 21536
rect 16114 21496 16120 21508
rect 16172 21496 16178 21548
rect 17129 21539 17187 21545
rect 17129 21505 17141 21539
rect 17175 21536 17187 21539
rect 17310 21536 17316 21548
rect 17175 21508 17316 21536
rect 17175 21505 17187 21508
rect 17129 21499 17187 21505
rect 17310 21496 17316 21508
rect 17368 21496 17374 21548
rect 17424 21539 17482 21545
rect 17424 21505 17436 21539
rect 17470 21534 17482 21539
rect 17604 21536 17632 21644
rect 18141 21641 18153 21675
rect 18187 21641 18199 21675
rect 20070 21672 20076 21684
rect 20031 21644 20076 21672
rect 18141 21635 18199 21641
rect 18156 21604 18184 21635
rect 20070 21632 20076 21644
rect 20128 21632 20134 21684
rect 22741 21675 22799 21681
rect 22741 21641 22753 21675
rect 22787 21672 22799 21675
rect 24026 21672 24032 21684
rect 22787 21644 24032 21672
rect 22787 21641 22799 21644
rect 22741 21635 22799 21641
rect 24026 21632 24032 21644
rect 24084 21632 24090 21684
rect 25406 21672 25412 21684
rect 24136 21644 25412 21672
rect 22186 21604 22192 21616
rect 18156 21576 22192 21604
rect 22186 21564 22192 21576
rect 22244 21564 22250 21616
rect 23382 21564 23388 21616
rect 23440 21564 23446 21616
rect 23658 21564 23664 21616
rect 23716 21604 23722 21616
rect 24136 21604 24164 21644
rect 25406 21632 25412 21644
rect 25464 21632 25470 21684
rect 27890 21672 27896 21684
rect 25884 21644 27896 21672
rect 23716 21576 24164 21604
rect 23716 21564 23722 21576
rect 18598 21536 18604 21548
rect 17512 21534 17632 21536
rect 17470 21508 17632 21534
rect 18559 21508 18604 21536
rect 17470 21506 17540 21508
rect 17470 21505 17482 21506
rect 17424 21499 17482 21505
rect 18598 21496 18604 21508
rect 18656 21496 18662 21548
rect 18874 21536 18880 21548
rect 18835 21508 18880 21536
rect 18874 21496 18880 21508
rect 18932 21496 18938 21548
rect 19334 21496 19340 21548
rect 19392 21536 19398 21548
rect 20257 21539 20315 21545
rect 20257 21536 20269 21539
rect 19392 21508 20269 21536
rect 19392 21496 19398 21508
rect 20257 21505 20269 21508
rect 20303 21505 20315 21539
rect 20257 21499 20315 21505
rect 20993 21539 21051 21545
rect 20993 21505 21005 21539
rect 21039 21536 21051 21539
rect 21818 21536 21824 21548
rect 21039 21508 21824 21536
rect 21039 21505 21051 21508
rect 20993 21499 21051 21505
rect 21818 21496 21824 21508
rect 21876 21496 21882 21548
rect 22554 21536 22560 21548
rect 22515 21508 22560 21536
rect 22554 21496 22560 21508
rect 22612 21496 22618 21548
rect 22833 21539 22891 21545
rect 22833 21505 22845 21539
rect 22879 21505 22891 21539
rect 22833 21499 22891 21505
rect 23293 21539 23351 21545
rect 23293 21505 23305 21539
rect 23339 21536 23351 21539
rect 23400 21536 23428 21564
rect 23339 21508 23428 21536
rect 23477 21539 23535 21545
rect 23339 21505 23351 21508
rect 23293 21499 23351 21505
rect 23477 21505 23489 21539
rect 23523 21536 23535 21539
rect 23566 21536 23572 21548
rect 23523 21508 23572 21536
rect 23523 21505 23535 21508
rect 23477 21499 23535 21505
rect 12802 21468 12808 21480
rect 12176 21440 12808 21468
rect 12802 21428 12808 21440
rect 12860 21428 12866 21480
rect 14918 21428 14924 21480
rect 14976 21468 14982 21480
rect 14976 21440 16712 21468
rect 14976 21428 14982 21440
rect 10134 21400 10140 21412
rect 8772 21372 10140 21400
rect 10134 21360 10140 21372
rect 10192 21360 10198 21412
rect 12342 21400 12348 21412
rect 12255 21372 12348 21400
rect 12342 21360 12348 21372
rect 12400 21360 12406 21412
rect 9858 21292 9864 21344
rect 9916 21332 9922 21344
rect 9953 21335 10011 21341
rect 9953 21332 9965 21335
rect 9916 21304 9965 21332
rect 9916 21292 9922 21304
rect 9953 21301 9965 21304
rect 9999 21301 10011 21335
rect 9953 21295 10011 21301
rect 11977 21335 12035 21341
rect 11977 21301 11989 21335
rect 12023 21332 12035 21335
rect 12250 21332 12256 21344
rect 12023 21304 12256 21332
rect 12023 21301 12035 21304
rect 11977 21295 12035 21301
rect 12250 21292 12256 21304
rect 12308 21292 12314 21344
rect 12360 21332 12388 21360
rect 14366 21332 14372 21344
rect 12360 21304 14372 21332
rect 14366 21292 14372 21304
rect 14424 21292 14430 21344
rect 15470 21292 15476 21344
rect 15528 21332 15534 21344
rect 15933 21335 15991 21341
rect 15933 21332 15945 21335
rect 15528 21304 15945 21332
rect 15528 21292 15534 21304
rect 15933 21301 15945 21304
rect 15979 21332 15991 21335
rect 16574 21332 16580 21344
rect 15979 21304 16580 21332
rect 15979 21301 15991 21304
rect 15933 21295 15991 21301
rect 16574 21292 16580 21304
rect 16632 21292 16638 21344
rect 16684 21332 16712 21440
rect 22848 21400 22876 21499
rect 23566 21496 23572 21508
rect 23624 21496 23630 21548
rect 24136 21545 24164 21576
rect 24394 21564 24400 21616
rect 24452 21604 24458 21616
rect 25777 21607 25835 21613
rect 25777 21604 25789 21607
rect 24452 21576 25789 21604
rect 24452 21564 24458 21576
rect 25777 21573 25789 21576
rect 25823 21573 25835 21607
rect 25777 21567 25835 21573
rect 24121 21539 24179 21545
rect 24121 21505 24133 21539
rect 24167 21505 24179 21539
rect 24121 21499 24179 21505
rect 24302 21496 24308 21548
rect 24360 21536 24366 21548
rect 24949 21539 25007 21545
rect 24360 21508 24405 21536
rect 24360 21496 24366 21508
rect 24949 21505 24961 21539
rect 24995 21505 25007 21539
rect 24949 21499 25007 21505
rect 25041 21539 25099 21545
rect 25041 21505 25053 21539
rect 25087 21505 25099 21539
rect 25222 21536 25228 21548
rect 25183 21508 25228 21536
rect 25041 21499 25099 21505
rect 23198 21400 23204 21412
rect 22848 21372 23204 21400
rect 23198 21360 23204 21372
rect 23256 21400 23262 21412
rect 24964 21400 24992 21499
rect 25056 21468 25084 21499
rect 25222 21496 25228 21508
rect 25280 21496 25286 21548
rect 25317 21539 25375 21545
rect 25317 21505 25329 21539
rect 25363 21536 25375 21539
rect 25884 21536 25912 21644
rect 27890 21632 27896 21644
rect 27948 21632 27954 21684
rect 27982 21632 27988 21684
rect 28040 21672 28046 21684
rect 28534 21672 28540 21684
rect 28040 21644 28540 21672
rect 28040 21632 28046 21644
rect 28534 21632 28540 21644
rect 28592 21632 28598 21684
rect 28626 21632 28632 21684
rect 28684 21672 28690 21684
rect 28905 21675 28963 21681
rect 28905 21672 28917 21675
rect 28684 21644 28917 21672
rect 28684 21632 28690 21644
rect 28905 21641 28917 21644
rect 28951 21641 28963 21675
rect 28905 21635 28963 21641
rect 28994 21632 29000 21684
rect 29052 21672 29058 21684
rect 29638 21672 29644 21684
rect 29052 21644 29644 21672
rect 29052 21632 29058 21644
rect 29638 21632 29644 21644
rect 29696 21632 29702 21684
rect 30006 21632 30012 21684
rect 30064 21672 30070 21684
rect 32490 21672 32496 21684
rect 30064 21644 32496 21672
rect 30064 21632 30070 21644
rect 32490 21632 32496 21644
rect 32548 21632 32554 21684
rect 34054 21672 34060 21684
rect 34015 21644 34060 21672
rect 34054 21632 34060 21644
rect 34112 21632 34118 21684
rect 37734 21632 37740 21684
rect 37792 21672 37798 21684
rect 37829 21675 37887 21681
rect 37829 21672 37841 21675
rect 37792 21644 37841 21672
rect 37792 21632 37798 21644
rect 37829 21641 37841 21644
rect 37875 21641 37887 21675
rect 37829 21635 37887 21641
rect 26418 21604 26424 21616
rect 26252 21576 26424 21604
rect 25363 21508 25912 21536
rect 25961 21539 26019 21545
rect 25363 21505 25375 21508
rect 25317 21499 25375 21505
rect 25961 21505 25973 21539
rect 26007 21505 26019 21539
rect 25961 21499 26019 21505
rect 25866 21468 25872 21480
rect 25056 21440 25872 21468
rect 25866 21428 25872 21440
rect 25924 21428 25930 21480
rect 25976 21468 26004 21499
rect 26050 21496 26056 21548
rect 26108 21536 26114 21548
rect 26252 21545 26280 21576
rect 26418 21564 26424 21576
rect 26476 21564 26482 21616
rect 27062 21564 27068 21616
rect 27120 21604 27126 21616
rect 27120 21576 28948 21604
rect 27120 21564 27126 21576
rect 28920 21548 28948 21576
rect 29086 21564 29092 21616
rect 29144 21604 29150 21616
rect 29914 21604 29920 21616
rect 29144 21576 29920 21604
rect 29144 21564 29150 21576
rect 26237 21539 26295 21545
rect 26108 21508 26153 21536
rect 26108 21496 26114 21508
rect 26237 21505 26249 21539
rect 26283 21505 26295 21539
rect 26237 21499 26295 21505
rect 26326 21496 26332 21548
rect 26384 21536 26390 21548
rect 26384 21508 26429 21536
rect 26384 21496 26390 21508
rect 27338 21496 27344 21548
rect 27396 21536 27402 21548
rect 27433 21539 27491 21545
rect 27433 21536 27445 21539
rect 27396 21508 27445 21536
rect 27396 21496 27402 21508
rect 27433 21505 27445 21508
rect 27479 21536 27491 21539
rect 28718 21536 28724 21548
rect 27479 21508 28724 21536
rect 27479 21505 27491 21508
rect 27433 21499 27491 21505
rect 28718 21496 28724 21508
rect 28776 21496 28782 21548
rect 28902 21496 28908 21548
rect 28960 21496 28966 21548
rect 28997 21539 29055 21545
rect 28997 21505 29009 21539
rect 29043 21536 29055 21539
rect 29178 21536 29184 21548
rect 29043 21508 29184 21536
rect 29043 21505 29055 21508
rect 28997 21499 29055 21505
rect 29178 21496 29184 21508
rect 29236 21496 29242 21548
rect 29362 21496 29368 21548
rect 29420 21536 29426 21548
rect 29748 21545 29776 21576
rect 29914 21564 29920 21576
rect 29972 21564 29978 21616
rect 31570 21604 31576 21616
rect 30944 21576 31576 21604
rect 30944 21548 30972 21576
rect 31570 21564 31576 21576
rect 31628 21604 31634 21616
rect 33689 21607 33747 21613
rect 31628 21576 32352 21604
rect 31628 21564 31634 21576
rect 29457 21539 29515 21545
rect 29457 21536 29469 21539
rect 29420 21508 29469 21536
rect 29420 21496 29426 21508
rect 29457 21505 29469 21508
rect 29503 21505 29515 21539
rect 29457 21499 29515 21505
rect 29733 21539 29791 21545
rect 29733 21505 29745 21539
rect 29779 21505 29791 21539
rect 29733 21499 29791 21505
rect 30837 21539 30895 21545
rect 30837 21505 30849 21539
rect 30883 21536 30895 21539
rect 30926 21536 30932 21548
rect 30883 21508 30932 21536
rect 30883 21505 30895 21508
rect 30837 21499 30895 21505
rect 30926 21496 30932 21508
rect 30984 21496 30990 21548
rect 31021 21539 31079 21545
rect 31021 21505 31033 21539
rect 31067 21505 31079 21539
rect 31021 21499 31079 21505
rect 31113 21539 31171 21545
rect 31113 21505 31125 21539
rect 31159 21536 31171 21539
rect 31294 21536 31300 21548
rect 31159 21508 31300 21536
rect 31159 21505 31171 21508
rect 31113 21499 31171 21505
rect 30558 21468 30564 21480
rect 25976 21440 27016 21468
rect 23256 21372 24992 21400
rect 23256 21360 23262 21372
rect 25222 21360 25228 21412
rect 25280 21400 25286 21412
rect 26326 21400 26332 21412
rect 25280 21372 26332 21400
rect 25280 21360 25286 21372
rect 26326 21360 26332 21372
rect 26384 21360 26390 21412
rect 26988 21400 27016 21440
rect 27453 21440 30564 21468
rect 27453 21400 27481 21440
rect 30558 21428 30564 21440
rect 30616 21428 30622 21480
rect 29546 21400 29552 21412
rect 26988 21372 27481 21400
rect 27724 21372 29552 21400
rect 19613 21335 19671 21341
rect 19613 21332 19625 21335
rect 16684 21304 19625 21332
rect 19613 21301 19625 21304
rect 19659 21301 19671 21335
rect 20806 21332 20812 21344
rect 20767 21304 20812 21332
rect 19613 21295 19671 21301
rect 20806 21292 20812 21304
rect 20864 21292 20870 21344
rect 22278 21292 22284 21344
rect 22336 21332 22342 21344
rect 22373 21335 22431 21341
rect 22373 21332 22385 21335
rect 22336 21304 22385 21332
rect 22336 21292 22342 21304
rect 22373 21301 22385 21304
rect 22419 21301 22431 21335
rect 22373 21295 22431 21301
rect 23106 21292 23112 21344
rect 23164 21332 23170 21344
rect 23661 21335 23719 21341
rect 23661 21332 23673 21335
rect 23164 21304 23673 21332
rect 23164 21292 23170 21304
rect 23661 21301 23673 21304
rect 23707 21301 23719 21335
rect 24118 21332 24124 21344
rect 24079 21304 24124 21332
rect 23661 21295 23719 21301
rect 24118 21292 24124 21304
rect 24176 21292 24182 21344
rect 24578 21292 24584 21344
rect 24636 21332 24642 21344
rect 24765 21335 24823 21341
rect 24765 21332 24777 21335
rect 24636 21304 24777 21332
rect 24636 21292 24642 21304
rect 24765 21301 24777 21304
rect 24811 21301 24823 21335
rect 24765 21295 24823 21301
rect 26050 21292 26056 21344
rect 26108 21332 26114 21344
rect 26234 21332 26240 21344
rect 26108 21304 26240 21332
rect 26108 21292 26114 21304
rect 26234 21292 26240 21304
rect 26292 21292 26298 21344
rect 27724 21341 27752 21372
rect 29546 21360 29552 21372
rect 29604 21360 29610 21412
rect 30742 21360 30748 21412
rect 30800 21400 30806 21412
rect 31036 21400 31064 21499
rect 31294 21496 31300 21508
rect 31352 21496 31358 21548
rect 32122 21536 32128 21548
rect 32083 21508 32128 21536
rect 32122 21496 32128 21508
rect 32180 21496 32186 21548
rect 32324 21545 32352 21576
rect 33689 21573 33701 21607
rect 33735 21604 33747 21607
rect 33962 21604 33968 21616
rect 33735 21576 33968 21604
rect 33735 21573 33747 21576
rect 33689 21567 33747 21573
rect 33962 21564 33968 21576
rect 34020 21564 34026 21616
rect 34517 21607 34575 21613
rect 34517 21573 34529 21607
rect 34563 21604 34575 21607
rect 34606 21604 34612 21616
rect 34563 21576 34612 21604
rect 34563 21573 34575 21576
rect 34517 21567 34575 21573
rect 34606 21564 34612 21576
rect 34664 21564 34670 21616
rect 34698 21564 34704 21616
rect 34756 21604 34762 21616
rect 34756 21576 36124 21604
rect 34756 21564 34762 21576
rect 36096 21548 36124 21576
rect 32309 21539 32367 21545
rect 32309 21505 32321 21539
rect 32355 21505 32367 21539
rect 32309 21499 32367 21505
rect 33873 21539 33931 21545
rect 33873 21505 33885 21539
rect 33919 21536 33931 21539
rect 34422 21536 34428 21548
rect 33919 21508 34428 21536
rect 33919 21505 33931 21508
rect 33873 21499 33931 21505
rect 34422 21496 34428 21508
rect 34480 21496 34486 21548
rect 35526 21496 35532 21548
rect 35584 21536 35590 21548
rect 35621 21539 35679 21545
rect 35621 21536 35633 21539
rect 35584 21508 35633 21536
rect 35584 21496 35590 21508
rect 35621 21505 35633 21508
rect 35667 21505 35679 21539
rect 35894 21536 35900 21548
rect 35855 21508 35900 21536
rect 35621 21499 35679 21505
rect 35894 21496 35900 21508
rect 35952 21496 35958 21548
rect 36078 21536 36084 21548
rect 36039 21508 36084 21536
rect 36078 21496 36084 21508
rect 36136 21496 36142 21548
rect 36357 21539 36415 21545
rect 36357 21505 36369 21539
rect 36403 21505 36415 21539
rect 36357 21499 36415 21505
rect 37461 21539 37519 21545
rect 37461 21505 37473 21539
rect 37507 21536 37519 21539
rect 37642 21536 37648 21548
rect 37507 21508 37648 21536
rect 37507 21505 37519 21508
rect 37461 21499 37519 21505
rect 34440 21468 34468 21496
rect 35710 21468 35716 21480
rect 34440 21440 35716 21468
rect 35710 21428 35716 21440
rect 35768 21468 35774 21480
rect 36372 21468 36400 21499
rect 37642 21496 37648 21508
rect 37700 21496 37706 21548
rect 37550 21468 37556 21480
rect 35768 21440 36400 21468
rect 37511 21440 37556 21468
rect 35768 21428 35774 21440
rect 37550 21428 37556 21440
rect 37608 21428 37614 21480
rect 31202 21400 31208 21412
rect 30800 21372 31208 21400
rect 30800 21360 30806 21372
rect 31202 21360 31208 21372
rect 31260 21360 31266 21412
rect 35986 21360 35992 21412
rect 36044 21400 36050 21412
rect 36173 21403 36231 21409
rect 36173 21400 36185 21403
rect 36044 21372 36185 21400
rect 36044 21360 36050 21372
rect 36173 21369 36185 21372
rect 36219 21369 36231 21403
rect 36173 21363 36231 21369
rect 27709 21335 27767 21341
rect 27709 21301 27721 21335
rect 27755 21301 27767 21335
rect 27890 21332 27896 21344
rect 27851 21304 27896 21332
rect 27709 21295 27767 21301
rect 27890 21292 27896 21304
rect 27948 21292 27954 21344
rect 28350 21292 28356 21344
rect 28408 21332 28414 21344
rect 28537 21335 28595 21341
rect 28537 21332 28549 21335
rect 28408 21304 28549 21332
rect 28408 21292 28414 21304
rect 28537 21301 28549 21304
rect 28583 21301 28595 21335
rect 28537 21295 28595 21301
rect 29457 21335 29515 21341
rect 29457 21301 29469 21335
rect 29503 21332 29515 21335
rect 29638 21332 29644 21344
rect 29503 21304 29644 21332
rect 29503 21301 29515 21304
rect 29457 21295 29515 21301
rect 29638 21292 29644 21304
rect 29696 21292 29702 21344
rect 30558 21292 30564 21344
rect 30616 21332 30622 21344
rect 30653 21335 30711 21341
rect 30653 21332 30665 21335
rect 30616 21304 30665 21332
rect 30616 21292 30622 21304
rect 30653 21301 30665 21304
rect 30699 21301 30711 21335
rect 30653 21295 30711 21301
rect 32125 21335 32183 21341
rect 32125 21301 32137 21335
rect 32171 21332 32183 21335
rect 32398 21332 32404 21344
rect 32171 21304 32404 21332
rect 32171 21301 32183 21304
rect 32125 21295 32183 21301
rect 32398 21292 32404 21304
rect 32456 21292 32462 21344
rect 34790 21292 34796 21344
rect 34848 21332 34854 21344
rect 34885 21335 34943 21341
rect 34885 21332 34897 21335
rect 34848 21304 34897 21332
rect 34848 21292 34854 21304
rect 34885 21301 34897 21304
rect 34931 21301 34943 21335
rect 34885 21295 34943 21301
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 9674 21128 9680 21140
rect 9416 21100 9680 21128
rect 8570 21060 8576 21072
rect 8128 21032 8576 21060
rect 8128 20933 8156 21032
rect 8570 21020 8576 21032
rect 8628 21020 8634 21072
rect 8389 20995 8447 21001
rect 8389 20961 8401 20995
rect 8435 20992 8447 20995
rect 9416 20992 9444 21100
rect 9674 21088 9680 21100
rect 9732 21088 9738 21140
rect 10134 21128 10140 21140
rect 10095 21100 10140 21128
rect 10134 21088 10140 21100
rect 10192 21088 10198 21140
rect 11790 21128 11796 21140
rect 11440 21100 11796 21128
rect 9493 21063 9551 21069
rect 9493 21029 9505 21063
rect 9539 21060 9551 21063
rect 9950 21060 9956 21072
rect 9539 21032 9956 21060
rect 9539 21029 9551 21032
rect 9493 21023 9551 21029
rect 9950 21020 9956 21032
rect 10008 21060 10014 21072
rect 10410 21060 10416 21072
rect 10008 21032 10416 21060
rect 10008 21020 10014 21032
rect 10410 21020 10416 21032
rect 10468 21020 10474 21072
rect 10594 21020 10600 21072
rect 10652 21020 10658 21072
rect 8435 20964 9444 20992
rect 9677 20995 9735 21001
rect 8435 20961 8447 20964
rect 8389 20955 8447 20961
rect 9677 20961 9689 20995
rect 9723 20992 9735 20995
rect 10042 20992 10048 21004
rect 9723 20964 10048 20992
rect 9723 20961 9735 20964
rect 9677 20955 9735 20961
rect 10042 20952 10048 20964
rect 10100 20952 10106 21004
rect 10226 20952 10232 21004
rect 10284 20992 10290 21004
rect 10612 20992 10640 21020
rect 11440 21001 11468 21100
rect 11790 21088 11796 21100
rect 11848 21128 11854 21140
rect 12802 21128 12808 21140
rect 11848 21100 12434 21128
rect 12763 21100 12808 21128
rect 11848 21088 11854 21100
rect 12406 21060 12434 21100
rect 12802 21088 12808 21100
rect 12860 21088 12866 21140
rect 13078 21088 13084 21140
rect 13136 21128 13142 21140
rect 13449 21131 13507 21137
rect 13449 21128 13461 21131
rect 13136 21100 13461 21128
rect 13136 21088 13142 21100
rect 13449 21097 13461 21100
rect 13495 21097 13507 21131
rect 13449 21091 13507 21097
rect 16482 21088 16488 21140
rect 16540 21128 16546 21140
rect 16669 21131 16727 21137
rect 16669 21128 16681 21131
rect 16540 21100 16681 21128
rect 16540 21088 16546 21100
rect 16669 21097 16681 21100
rect 16715 21128 16727 21131
rect 16942 21128 16948 21140
rect 16715 21100 16948 21128
rect 16715 21097 16727 21100
rect 16669 21091 16727 21097
rect 16942 21088 16948 21100
rect 17000 21088 17006 21140
rect 19245 21131 19303 21137
rect 19245 21128 19257 21131
rect 17696 21100 19257 21128
rect 13170 21060 13176 21072
rect 12406 21032 13176 21060
rect 13170 21020 13176 21032
rect 13228 21020 13234 21072
rect 15654 21020 15660 21072
rect 15712 21060 15718 21072
rect 16206 21060 16212 21072
rect 15712 21032 16212 21060
rect 15712 21020 15718 21032
rect 16206 21020 16212 21032
rect 16264 21060 16270 21072
rect 16301 21063 16359 21069
rect 16301 21060 16313 21063
rect 16264 21032 16313 21060
rect 16264 21020 16270 21032
rect 16301 21029 16313 21032
rect 16347 21029 16359 21063
rect 16301 21023 16359 21029
rect 11425 20995 11483 21001
rect 10284 20964 10456 20992
rect 10612 20964 10824 20992
rect 10284 20952 10290 20964
rect 8113 20927 8171 20933
rect 8113 20893 8125 20927
rect 8159 20893 8171 20927
rect 8113 20887 8171 20893
rect 8205 20927 8263 20933
rect 8205 20893 8217 20927
rect 8251 20893 8263 20927
rect 8205 20887 8263 20893
rect 9401 20927 9459 20933
rect 9401 20893 9413 20927
rect 9447 20924 9459 20927
rect 9766 20924 9772 20936
rect 9447 20896 9772 20924
rect 9447 20893 9459 20896
rect 9401 20887 9459 20893
rect 8220 20856 8248 20887
rect 9766 20884 9772 20896
rect 9824 20924 9830 20936
rect 10318 20924 10324 20936
rect 9824 20896 10324 20924
rect 9824 20884 9830 20896
rect 10318 20884 10324 20896
rect 10376 20884 10382 20936
rect 10428 20933 10456 20964
rect 10413 20927 10471 20933
rect 10413 20893 10425 20927
rect 10459 20893 10471 20927
rect 10413 20887 10471 20893
rect 10505 20927 10563 20933
rect 10505 20893 10517 20927
rect 10551 20893 10563 20927
rect 10505 20887 10563 20893
rect 9858 20856 9864 20868
rect 8220 20828 9864 20856
rect 9858 20816 9864 20828
rect 9916 20816 9922 20868
rect 10520 20856 10548 20887
rect 10594 20884 10600 20936
rect 10652 20924 10658 20936
rect 10796 20933 10824 20964
rect 11425 20961 11437 20995
rect 11471 20961 11483 20995
rect 11425 20955 11483 20961
rect 13354 20952 13360 21004
rect 13412 20992 13418 21004
rect 13412 20964 14596 20992
rect 13412 20952 13418 20964
rect 10781 20927 10839 20933
rect 10652 20896 10697 20924
rect 10652 20884 10658 20896
rect 10781 20893 10793 20927
rect 10827 20924 10839 20927
rect 11330 20924 11336 20936
rect 10827 20896 11336 20924
rect 10827 20893 10839 20896
rect 10781 20887 10839 20893
rect 11330 20884 11336 20896
rect 11388 20884 11394 20936
rect 11698 20933 11704 20936
rect 11692 20924 11704 20933
rect 11659 20896 11704 20924
rect 11692 20887 11704 20896
rect 11698 20884 11704 20887
rect 11756 20884 11762 20936
rect 14366 20884 14372 20936
rect 14424 20924 14430 20936
rect 14461 20927 14519 20933
rect 14461 20924 14473 20927
rect 14424 20896 14473 20924
rect 14424 20884 14430 20896
rect 14461 20893 14473 20896
rect 14507 20893 14519 20927
rect 14568 20924 14596 20964
rect 17310 20952 17316 21004
rect 17368 20992 17374 21004
rect 17696 21001 17724 21100
rect 19245 21097 19257 21100
rect 19291 21097 19303 21131
rect 19245 21091 19303 21097
rect 22554 21088 22560 21140
rect 22612 21128 22618 21140
rect 27614 21128 27620 21140
rect 22612 21100 27620 21128
rect 22612 21088 22618 21100
rect 27614 21088 27620 21100
rect 27672 21088 27678 21140
rect 27706 21088 27712 21140
rect 27764 21128 27770 21140
rect 30009 21131 30067 21137
rect 30009 21128 30021 21131
rect 27764 21100 30021 21128
rect 27764 21088 27770 21100
rect 30009 21097 30021 21100
rect 30055 21097 30067 21131
rect 33318 21128 33324 21140
rect 30009 21091 30067 21097
rect 30760 21100 33180 21128
rect 33279 21100 33324 21128
rect 22186 21020 22192 21072
rect 22244 21060 22250 21072
rect 23658 21060 23664 21072
rect 22244 21032 23664 21060
rect 22244 21020 22250 21032
rect 23658 21020 23664 21032
rect 23716 21020 23722 21072
rect 30561 21063 30619 21069
rect 30561 21060 30573 21063
rect 23768 21032 28028 21060
rect 17681 20995 17739 21001
rect 17681 20992 17693 20995
rect 17368 20964 17693 20992
rect 17368 20952 17374 20964
rect 17681 20961 17693 20964
rect 17727 20961 17739 20995
rect 17681 20955 17739 20961
rect 21634 20952 21640 21004
rect 21692 20992 21698 21004
rect 21821 20995 21879 21001
rect 21821 20992 21833 20995
rect 21692 20964 21833 20992
rect 21692 20952 21698 20964
rect 21821 20961 21833 20964
rect 21867 20961 21879 20995
rect 22462 20992 22468 21004
rect 21821 20955 21879 20961
rect 22112 20964 22468 20992
rect 14717 20927 14775 20933
rect 14717 20924 14729 20927
rect 14568 20896 14729 20924
rect 14461 20887 14519 20893
rect 14717 20893 14729 20896
rect 14763 20893 14775 20927
rect 17957 20927 18015 20933
rect 17957 20924 17969 20927
rect 14717 20887 14775 20893
rect 14844 20896 17969 20924
rect 11974 20856 11980 20868
rect 10520 20828 11980 20856
rect 11974 20816 11980 20828
rect 12032 20816 12038 20868
rect 12802 20816 12808 20868
rect 12860 20856 12866 20868
rect 13357 20859 13415 20865
rect 13357 20856 13369 20859
rect 12860 20828 13369 20856
rect 12860 20816 12866 20828
rect 13357 20825 13369 20828
rect 13403 20825 13415 20859
rect 13357 20819 13415 20825
rect 13446 20816 13452 20868
rect 13504 20856 13510 20868
rect 14844 20856 14872 20896
rect 17957 20893 17969 20896
rect 18003 20893 18015 20927
rect 17957 20887 18015 20893
rect 19429 20927 19487 20933
rect 19429 20893 19441 20927
rect 19475 20893 19487 20927
rect 19429 20887 19487 20893
rect 19889 20927 19947 20933
rect 19889 20893 19901 20927
rect 19935 20924 19947 20927
rect 20070 20924 20076 20936
rect 19935 20896 20076 20924
rect 19935 20893 19947 20896
rect 19889 20887 19947 20893
rect 19444 20856 19472 20887
rect 20070 20884 20076 20896
rect 20128 20884 20134 20936
rect 20165 20927 20223 20933
rect 20165 20893 20177 20927
rect 20211 20924 20223 20927
rect 21726 20924 21732 20936
rect 20211 20896 21732 20924
rect 20211 20893 20223 20896
rect 20165 20887 20223 20893
rect 21726 20884 21732 20896
rect 21784 20884 21790 20936
rect 22112 20933 22140 20964
rect 22462 20952 22468 20964
rect 22520 20992 22526 21004
rect 22520 20964 23612 20992
rect 22520 20952 22526 20964
rect 23584 20936 23612 20964
rect 22097 20927 22155 20933
rect 22097 20893 22109 20927
rect 22143 20893 22155 20927
rect 22097 20887 22155 20893
rect 23106 20884 23112 20936
rect 23164 20924 23170 20936
rect 23339 20927 23397 20933
rect 23339 20924 23351 20927
rect 23164 20896 23351 20924
rect 23164 20884 23170 20896
rect 23339 20893 23351 20896
rect 23385 20893 23397 20927
rect 23471 20921 23477 20933
rect 23432 20893 23477 20921
rect 23339 20887 23397 20893
rect 23471 20881 23477 20893
rect 23529 20881 23535 20933
rect 23566 20884 23572 20936
rect 23624 20924 23630 20936
rect 23768 20933 23796 21032
rect 24118 20952 24124 21004
rect 24176 20992 24182 21004
rect 24765 20995 24823 21001
rect 24765 20992 24777 20995
rect 24176 20964 24777 20992
rect 24176 20952 24182 20964
rect 24765 20961 24777 20964
rect 24811 20992 24823 20995
rect 24946 20992 24952 21004
rect 24811 20964 24952 20992
rect 24811 20961 24823 20964
rect 24765 20955 24823 20961
rect 24946 20952 24952 20964
rect 25004 20952 25010 21004
rect 25041 20995 25099 21001
rect 25041 20961 25053 20995
rect 25087 20992 25099 20995
rect 25222 20992 25228 21004
rect 25087 20964 25228 20992
rect 25087 20961 25099 20964
rect 25041 20955 25099 20961
rect 25222 20952 25228 20964
rect 25280 20952 25286 21004
rect 26326 20952 26332 21004
rect 26384 20992 26390 21004
rect 26881 20995 26939 21001
rect 26881 20992 26893 20995
rect 26384 20964 26893 20992
rect 26384 20952 26390 20964
rect 26881 20961 26893 20964
rect 26927 20992 26939 20995
rect 27062 20992 27068 21004
rect 26927 20964 27068 20992
rect 26927 20961 26939 20964
rect 26881 20955 26939 20961
rect 27062 20952 27068 20964
rect 27120 20952 27126 21004
rect 27341 20995 27399 21001
rect 27341 20961 27353 20995
rect 27387 20992 27399 20995
rect 27890 20992 27896 21004
rect 27387 20964 27896 20992
rect 27387 20961 27399 20964
rect 27341 20955 27399 20961
rect 27890 20952 27896 20964
rect 27948 20952 27954 21004
rect 28000 20992 28028 21032
rect 28184 21032 30573 21060
rect 28184 20992 28212 21032
rect 30561 21029 30573 21032
rect 30607 21029 30619 21063
rect 30561 21023 30619 21029
rect 28000 20964 28212 20992
rect 28442 20952 28448 21004
rect 28500 20992 28506 21004
rect 29638 20992 29644 21004
rect 28500 20964 29224 20992
rect 29599 20964 29644 20992
rect 28500 20952 28506 20964
rect 23753 20927 23811 20933
rect 23624 20896 23669 20924
rect 23624 20884 23630 20896
rect 23753 20893 23765 20927
rect 23799 20893 23811 20927
rect 23753 20887 23811 20893
rect 26237 20927 26295 20933
rect 26237 20893 26249 20927
rect 26283 20924 26295 20927
rect 26786 20924 26792 20936
rect 26283 20896 26792 20924
rect 26283 20893 26295 20896
rect 26237 20887 26295 20893
rect 26786 20884 26792 20896
rect 26844 20884 26850 20936
rect 27249 20927 27307 20933
rect 27249 20893 27261 20927
rect 27295 20924 27307 20927
rect 27295 20921 28212 20924
rect 28350 20921 28356 20936
rect 27295 20896 28356 20921
rect 27295 20893 27307 20896
rect 28184 20893 28356 20896
rect 28408 20924 28414 20936
rect 28408 20896 28453 20924
rect 27249 20887 27307 20893
rect 28350 20884 28356 20893
rect 28408 20884 28414 20896
rect 28534 20884 28540 20936
rect 28592 20924 28598 20936
rect 28813 20927 28871 20933
rect 28813 20924 28825 20927
rect 28592 20896 28825 20924
rect 28592 20884 28598 20896
rect 28813 20893 28825 20896
rect 28859 20893 28871 20927
rect 28813 20887 28871 20893
rect 28902 20884 28908 20936
rect 28960 20924 28966 20936
rect 28997 20927 29055 20933
rect 28997 20924 29009 20927
rect 28960 20896 29009 20924
rect 28960 20884 28966 20896
rect 28997 20893 29009 20896
rect 29043 20893 29055 20927
rect 28997 20887 29055 20893
rect 13504 20828 14872 20856
rect 16868 20828 19472 20856
rect 13504 20816 13510 20828
rect 8386 20788 8392 20800
rect 8347 20760 8392 20788
rect 8386 20748 8392 20760
rect 8444 20748 8450 20800
rect 9674 20788 9680 20800
rect 9635 20760 9680 20788
rect 9674 20748 9680 20760
rect 9732 20748 9738 20800
rect 9766 20748 9772 20800
rect 9824 20788 9830 20800
rect 10962 20788 10968 20800
rect 9824 20760 10968 20788
rect 9824 20748 9830 20760
rect 10962 20748 10968 20760
rect 11020 20788 11026 20800
rect 12618 20788 12624 20800
rect 11020 20760 12624 20788
rect 11020 20748 11026 20760
rect 12618 20748 12624 20760
rect 12676 20748 12682 20800
rect 13630 20748 13636 20800
rect 13688 20788 13694 20800
rect 14274 20788 14280 20800
rect 13688 20760 14280 20788
rect 13688 20748 13694 20760
rect 14274 20748 14280 20760
rect 14332 20748 14338 20800
rect 15841 20791 15899 20797
rect 15841 20757 15853 20791
rect 15887 20788 15899 20791
rect 15930 20788 15936 20800
rect 15887 20760 15936 20788
rect 15887 20757 15899 20760
rect 15841 20751 15899 20757
rect 15930 20748 15936 20760
rect 15988 20788 15994 20800
rect 16868 20797 16896 20828
rect 27890 20816 27896 20868
rect 27948 20856 27954 20868
rect 27948 20828 28028 20856
rect 27948 20816 27954 20828
rect 16669 20791 16727 20797
rect 16669 20788 16681 20791
rect 15988 20760 16681 20788
rect 15988 20748 15994 20760
rect 16669 20757 16681 20760
rect 16715 20757 16727 20791
rect 16669 20751 16727 20757
rect 16853 20791 16911 20797
rect 16853 20757 16865 20791
rect 16899 20757 16911 20791
rect 16853 20751 16911 20757
rect 18693 20791 18751 20797
rect 18693 20757 18705 20791
rect 18739 20788 18751 20791
rect 20714 20788 20720 20800
rect 18739 20760 20720 20788
rect 18739 20757 18751 20760
rect 18693 20751 18751 20757
rect 20714 20748 20720 20760
rect 20772 20748 20778 20800
rect 20898 20788 20904 20800
rect 20859 20760 20904 20788
rect 20898 20748 20904 20760
rect 20956 20748 20962 20800
rect 23106 20788 23112 20800
rect 23067 20760 23112 20788
rect 23106 20748 23112 20760
rect 23164 20748 23170 20800
rect 24854 20748 24860 20800
rect 24912 20788 24918 20800
rect 25590 20788 25596 20800
rect 24912 20760 25596 20788
rect 24912 20748 24918 20760
rect 25590 20748 25596 20760
rect 25648 20788 25654 20800
rect 26329 20791 26387 20797
rect 26329 20788 26341 20791
rect 25648 20760 26341 20788
rect 25648 20748 25654 20760
rect 26329 20757 26341 20760
rect 26375 20757 26387 20791
rect 26329 20751 26387 20757
rect 26418 20748 26424 20800
rect 26476 20788 26482 20800
rect 27525 20791 27583 20797
rect 27525 20788 27537 20791
rect 26476 20760 27537 20788
rect 26476 20748 26482 20760
rect 27525 20757 27537 20760
rect 27571 20757 27583 20791
rect 28000 20788 28028 20828
rect 28074 20816 28080 20868
rect 28132 20856 28138 20868
rect 28261 20859 28319 20865
rect 28132 20828 28177 20856
rect 28132 20816 28138 20828
rect 28261 20825 28273 20859
rect 28307 20856 28319 20859
rect 28442 20856 28448 20868
rect 28307 20828 28448 20856
rect 28307 20825 28319 20828
rect 28261 20819 28319 20825
rect 28442 20816 28448 20828
rect 28500 20816 28506 20868
rect 29196 20856 29224 20964
rect 29638 20952 29644 20964
rect 29696 20952 29702 21004
rect 30760 21001 30788 21100
rect 33042 21060 33048 21072
rect 30852 21032 33048 21060
rect 30852 21001 30880 21032
rect 33042 21020 33048 21032
rect 33100 21020 33106 21072
rect 33152 21060 33180 21100
rect 33318 21088 33324 21100
rect 33376 21088 33382 21140
rect 37001 21131 37059 21137
rect 37001 21128 37013 21131
rect 34992 21100 37013 21128
rect 34882 21060 34888 21072
rect 33152 21032 34888 21060
rect 34882 21020 34888 21032
rect 34940 21020 34946 21072
rect 30745 20995 30803 21001
rect 30745 20961 30757 20995
rect 30791 20961 30803 20995
rect 30745 20955 30803 20961
rect 30837 20995 30895 21001
rect 30837 20961 30849 20995
rect 30883 20961 30895 20995
rect 31018 20992 31024 21004
rect 30979 20964 31024 20992
rect 30837 20955 30895 20961
rect 31018 20952 31024 20964
rect 31076 20952 31082 21004
rect 31570 20992 31576 21004
rect 31531 20964 31576 20992
rect 31570 20952 31576 20964
rect 31628 20952 31634 21004
rect 34606 20952 34612 21004
rect 34664 20992 34670 21004
rect 34992 21001 35020 21100
rect 37001 21097 37013 21100
rect 37047 21097 37059 21131
rect 37642 21128 37648 21140
rect 37603 21100 37648 21128
rect 37001 21091 37059 21097
rect 37642 21088 37648 21100
rect 37700 21088 37706 21140
rect 35618 21020 35624 21072
rect 35676 21020 35682 21072
rect 35894 21020 35900 21072
rect 35952 21020 35958 21072
rect 35986 21020 35992 21072
rect 36044 21060 36050 21072
rect 37553 21063 37611 21069
rect 37553 21060 37565 21063
rect 36044 21032 36676 21060
rect 36044 21020 36050 21032
rect 34977 20995 35035 21001
rect 34977 20992 34989 20995
rect 34664 20964 34989 20992
rect 34664 20952 34670 20964
rect 34977 20961 34989 20964
rect 35023 20961 35035 20995
rect 35636 20992 35664 21020
rect 35912 20992 35940 21020
rect 34977 20955 35035 20961
rect 35084 20964 35664 20992
rect 35728 20964 35940 20992
rect 29270 20884 29276 20936
rect 29328 20924 29334 20936
rect 29733 20927 29791 20933
rect 29733 20924 29745 20927
rect 29328 20896 29745 20924
rect 29328 20884 29334 20896
rect 29733 20893 29745 20896
rect 29779 20893 29791 20927
rect 30926 20924 30932 20936
rect 30887 20896 30932 20924
rect 29733 20887 29791 20893
rect 30926 20884 30932 20896
rect 30984 20884 30990 20936
rect 31757 20927 31815 20933
rect 31757 20893 31769 20927
rect 31803 20924 31815 20927
rect 32122 20924 32128 20936
rect 31803 20896 32128 20924
rect 31803 20893 31815 20896
rect 31757 20887 31815 20893
rect 32122 20884 32128 20896
rect 32180 20884 32186 20936
rect 32398 20924 32404 20936
rect 32359 20896 32404 20924
rect 32398 20884 32404 20896
rect 32456 20884 32462 20936
rect 33226 20924 33232 20936
rect 33187 20896 33232 20924
rect 33226 20884 33232 20896
rect 33284 20884 33290 20936
rect 33321 20927 33379 20933
rect 33321 20893 33333 20927
rect 33367 20893 33379 20927
rect 34698 20924 34704 20936
rect 34659 20896 34704 20924
rect 33321 20887 33379 20893
rect 30742 20856 30748 20868
rect 29196 20828 30748 20856
rect 30742 20816 30748 20828
rect 30800 20816 30806 20868
rect 31941 20859 31999 20865
rect 31941 20825 31953 20859
rect 31987 20856 31999 20859
rect 32490 20856 32496 20868
rect 31987 20828 32496 20856
rect 31987 20825 31999 20828
rect 31941 20819 31999 20825
rect 32490 20816 32496 20828
rect 32548 20856 32554 20868
rect 32585 20859 32643 20865
rect 32585 20856 32597 20859
rect 32548 20828 32597 20856
rect 32548 20816 32554 20828
rect 32585 20825 32597 20828
rect 32631 20856 32643 20859
rect 33336 20856 33364 20887
rect 34698 20884 34704 20896
rect 34756 20884 34762 20936
rect 34793 20927 34851 20933
rect 34793 20893 34805 20927
rect 34839 20924 34851 20927
rect 35084 20924 35112 20964
rect 34839 20896 35112 20924
rect 34839 20893 34851 20896
rect 34793 20887 34851 20893
rect 35526 20884 35532 20936
rect 35584 20924 35590 20936
rect 35728 20933 35756 20964
rect 35621 20927 35679 20933
rect 35621 20924 35633 20927
rect 35584 20896 35633 20924
rect 35584 20884 35590 20896
rect 35621 20893 35633 20896
rect 35667 20893 35679 20927
rect 35621 20887 35679 20893
rect 35713 20927 35771 20933
rect 35713 20893 35725 20927
rect 35759 20893 35771 20927
rect 35894 20924 35900 20936
rect 35855 20896 35900 20924
rect 35713 20887 35771 20893
rect 35894 20884 35900 20896
rect 35952 20884 35958 20936
rect 35989 20927 36047 20933
rect 35989 20893 36001 20927
rect 36035 20924 36047 20927
rect 36078 20924 36084 20936
rect 36035 20896 36084 20924
rect 36035 20893 36047 20896
rect 35989 20887 36047 20893
rect 36078 20884 36084 20896
rect 36136 20884 36142 20936
rect 36648 20933 36676 21032
rect 36740 21032 37565 21060
rect 36740 21001 36768 21032
rect 37553 21029 37565 21032
rect 37599 21060 37611 21063
rect 37826 21060 37832 21072
rect 37599 21032 37832 21060
rect 37599 21029 37611 21032
rect 37553 21023 37611 21029
rect 37826 21020 37832 21032
rect 37884 21020 37890 21072
rect 36725 20995 36783 21001
rect 36725 20961 36737 20995
rect 36771 20961 36783 20995
rect 37737 20995 37795 21001
rect 37737 20992 37749 20995
rect 36725 20955 36783 20961
rect 37568 20964 37749 20992
rect 36633 20927 36691 20933
rect 36633 20893 36645 20927
rect 36679 20924 36691 20927
rect 37461 20927 37519 20933
rect 37461 20924 37473 20927
rect 36679 20896 37473 20924
rect 36679 20893 36691 20896
rect 36633 20887 36691 20893
rect 37461 20893 37473 20896
rect 37507 20893 37519 20927
rect 37461 20887 37519 20893
rect 32631 20828 33364 20856
rect 32631 20825 32643 20828
rect 32585 20819 32643 20825
rect 34882 20816 34888 20868
rect 34940 20856 34946 20868
rect 37568 20856 37596 20964
rect 37737 20961 37749 20964
rect 37783 20961 37795 20995
rect 37737 20955 37795 20961
rect 34940 20828 37596 20856
rect 34940 20816 34946 20828
rect 28175 20791 28233 20797
rect 28175 20788 28187 20791
rect 28000 20760 28187 20788
rect 27525 20751 27583 20757
rect 28175 20757 28187 20760
rect 28221 20757 28233 20791
rect 28175 20751 28233 20757
rect 28905 20791 28963 20797
rect 28905 20757 28917 20791
rect 28951 20788 28963 20791
rect 29178 20788 29184 20800
rect 28951 20760 29184 20788
rect 28951 20757 28963 20760
rect 28905 20751 28963 20757
rect 29178 20748 29184 20760
rect 29236 20748 29242 20800
rect 29362 20748 29368 20800
rect 29420 20788 29426 20800
rect 31662 20788 31668 20800
rect 29420 20760 31668 20788
rect 29420 20748 29426 20760
rect 31662 20748 31668 20760
rect 31720 20748 31726 20800
rect 32030 20748 32036 20800
rect 32088 20788 32094 20800
rect 32769 20791 32827 20797
rect 32769 20788 32781 20791
rect 32088 20760 32781 20788
rect 32088 20748 32094 20760
rect 32769 20757 32781 20760
rect 32815 20757 32827 20791
rect 32769 20751 32827 20757
rect 33134 20748 33140 20800
rect 33192 20788 33198 20800
rect 33597 20791 33655 20797
rect 33597 20788 33609 20791
rect 33192 20760 33609 20788
rect 33192 20748 33198 20760
rect 33597 20757 33609 20760
rect 33643 20757 33655 20791
rect 35434 20788 35440 20800
rect 35395 20760 35440 20788
rect 33597 20751 33655 20757
rect 35434 20748 35440 20760
rect 35492 20748 35498 20800
rect 35710 20748 35716 20800
rect 35768 20788 35774 20800
rect 35894 20788 35900 20800
rect 35768 20760 35900 20788
rect 35768 20748 35774 20760
rect 35894 20748 35900 20760
rect 35952 20748 35958 20800
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 9953 20587 10011 20593
rect 9953 20553 9965 20587
rect 9999 20584 10011 20587
rect 10594 20584 10600 20596
rect 9999 20556 10600 20584
rect 9999 20553 10011 20556
rect 9953 20547 10011 20553
rect 10594 20544 10600 20556
rect 10652 20544 10658 20596
rect 13173 20587 13231 20593
rect 13173 20553 13185 20587
rect 13219 20584 13231 20587
rect 13262 20584 13268 20596
rect 13219 20556 13268 20584
rect 13219 20553 13231 20556
rect 13173 20547 13231 20553
rect 13262 20544 13268 20556
rect 13320 20544 13326 20596
rect 14090 20544 14096 20596
rect 14148 20584 14154 20596
rect 14829 20587 14887 20593
rect 14829 20584 14841 20587
rect 14148 20556 14841 20584
rect 14148 20544 14154 20556
rect 14829 20553 14841 20556
rect 14875 20553 14887 20587
rect 15286 20584 15292 20596
rect 15247 20556 15292 20584
rect 14829 20547 14887 20553
rect 15286 20544 15292 20556
rect 15344 20544 15350 20596
rect 17310 20584 17316 20596
rect 17271 20556 17316 20584
rect 17310 20544 17316 20556
rect 17368 20544 17374 20596
rect 19245 20587 19303 20593
rect 19245 20553 19257 20587
rect 19291 20584 19303 20587
rect 19426 20584 19432 20596
rect 19291 20556 19432 20584
rect 19291 20553 19303 20556
rect 19245 20547 19303 20553
rect 19426 20544 19432 20556
rect 19484 20544 19490 20596
rect 20990 20584 20996 20596
rect 20088 20556 20996 20584
rect 20088 20528 20116 20556
rect 20990 20544 20996 20556
rect 21048 20544 21054 20596
rect 21726 20544 21732 20596
rect 21784 20584 21790 20596
rect 21821 20587 21879 20593
rect 21821 20584 21833 20587
rect 21784 20556 21833 20584
rect 21784 20544 21790 20556
rect 21821 20553 21833 20556
rect 21867 20553 21879 20587
rect 21821 20547 21879 20553
rect 21910 20544 21916 20596
rect 21968 20584 21974 20596
rect 22925 20587 22983 20593
rect 22925 20584 22937 20587
rect 21968 20556 22937 20584
rect 21968 20544 21974 20556
rect 22925 20553 22937 20556
rect 22971 20553 22983 20587
rect 22925 20547 22983 20553
rect 23566 20544 23572 20596
rect 23624 20584 23630 20596
rect 23624 20556 25636 20584
rect 23624 20544 23630 20556
rect 10042 20516 10048 20528
rect 9048 20488 10048 20516
rect 8386 20408 8392 20460
rect 8444 20448 8450 20460
rect 8665 20451 8723 20457
rect 8665 20448 8677 20451
rect 8444 20420 8677 20448
rect 8444 20408 8450 20420
rect 8665 20417 8677 20420
rect 8711 20417 8723 20451
rect 9048 20448 9076 20488
rect 10042 20476 10048 20488
rect 10100 20476 10106 20528
rect 17221 20519 17279 20525
rect 11900 20488 14412 20516
rect 8665 20411 8723 20417
rect 8864 20420 9076 20448
rect 7561 20383 7619 20389
rect 7561 20349 7573 20383
rect 7607 20380 7619 20383
rect 7742 20380 7748 20392
rect 7607 20352 7748 20380
rect 7607 20349 7619 20352
rect 7561 20343 7619 20349
rect 7742 20340 7748 20352
rect 7800 20340 7806 20392
rect 8754 20380 8760 20392
rect 8715 20352 8760 20380
rect 8754 20340 8760 20352
rect 8812 20340 8818 20392
rect 8864 20389 8892 20420
rect 9674 20408 9680 20460
rect 9732 20448 9738 20460
rect 10137 20451 10195 20457
rect 10137 20448 10149 20451
rect 9732 20420 10149 20448
rect 9732 20408 9738 20420
rect 10137 20417 10149 20420
rect 10183 20417 10195 20451
rect 10318 20448 10324 20460
rect 10279 20420 10324 20448
rect 10137 20411 10195 20417
rect 10318 20408 10324 20420
rect 10376 20408 10382 20460
rect 10410 20408 10416 20460
rect 10468 20448 10474 20460
rect 10468 20420 10513 20448
rect 10468 20408 10474 20420
rect 10962 20408 10968 20460
rect 11020 20448 11026 20460
rect 11900 20457 11928 20488
rect 11885 20451 11943 20457
rect 11885 20448 11897 20451
rect 11020 20420 11897 20448
rect 11020 20408 11026 20420
rect 11885 20417 11897 20420
rect 11931 20417 11943 20451
rect 11885 20411 11943 20417
rect 13357 20451 13415 20457
rect 13357 20417 13369 20451
rect 13403 20448 13415 20451
rect 14093 20451 14151 20457
rect 13403 20420 13860 20448
rect 13403 20417 13415 20420
rect 13357 20411 13415 20417
rect 8849 20383 8907 20389
rect 8849 20349 8861 20383
rect 8895 20349 8907 20383
rect 8849 20343 8907 20349
rect 8941 20383 8999 20389
rect 8941 20349 8953 20383
rect 8987 20349 8999 20383
rect 12158 20380 12164 20392
rect 12119 20352 12164 20380
rect 8941 20343 8999 20349
rect 7929 20315 7987 20321
rect 7929 20281 7941 20315
rect 7975 20312 7987 20315
rect 8481 20315 8539 20321
rect 8481 20312 8493 20315
rect 7975 20284 8493 20312
rect 7975 20281 7987 20284
rect 7929 20275 7987 20281
rect 8481 20281 8493 20284
rect 8527 20281 8539 20315
rect 8481 20275 8539 20281
rect 8021 20247 8079 20253
rect 8021 20213 8033 20247
rect 8067 20244 8079 20247
rect 8294 20244 8300 20256
rect 8067 20216 8300 20244
rect 8067 20213 8079 20216
rect 8021 20207 8079 20213
rect 8294 20204 8300 20216
rect 8352 20204 8358 20256
rect 8956 20244 8984 20343
rect 12158 20340 12164 20352
rect 12216 20340 12222 20392
rect 13630 20340 13636 20392
rect 13688 20380 13694 20392
rect 13688 20352 13733 20380
rect 13688 20340 13694 20352
rect 11974 20272 11980 20324
rect 12032 20312 12038 20324
rect 13541 20315 13599 20321
rect 13541 20312 13553 20315
rect 12032 20284 13553 20312
rect 12032 20272 12038 20284
rect 13541 20281 13553 20284
rect 13587 20281 13599 20315
rect 13832 20312 13860 20420
rect 14093 20417 14105 20451
rect 14139 20417 14151 20451
rect 14274 20448 14280 20460
rect 14235 20420 14280 20448
rect 14093 20411 14151 20417
rect 14108 20380 14136 20411
rect 14274 20408 14280 20420
rect 14332 20408 14338 20460
rect 14384 20457 14412 20488
rect 17221 20485 17233 20519
rect 17267 20516 17279 20519
rect 17862 20516 17868 20528
rect 17267 20488 17868 20516
rect 17267 20485 17279 20488
rect 17221 20479 17279 20485
rect 17862 20476 17868 20488
rect 17920 20516 17926 20528
rect 18417 20519 18475 20525
rect 18417 20516 18429 20519
rect 17920 20488 18429 20516
rect 17920 20476 17926 20488
rect 18417 20485 18429 20488
rect 18463 20485 18475 20519
rect 18417 20479 18475 20485
rect 18690 20476 18696 20528
rect 18748 20516 18754 20528
rect 18877 20519 18935 20525
rect 18877 20516 18889 20519
rect 18748 20488 18889 20516
rect 18748 20476 18754 20488
rect 18877 20485 18889 20488
rect 18923 20485 18935 20519
rect 18877 20479 18935 20485
rect 18966 20476 18972 20528
rect 19024 20516 19030 20528
rect 19077 20519 19135 20525
rect 19077 20516 19089 20519
rect 19024 20488 19089 20516
rect 19024 20476 19030 20488
rect 19077 20485 19089 20488
rect 19123 20485 19135 20519
rect 19077 20479 19135 20485
rect 20070 20476 20076 20528
rect 20128 20476 20134 20528
rect 20714 20476 20720 20528
rect 20772 20516 20778 20528
rect 20772 20488 21128 20516
rect 20772 20476 20778 20488
rect 14369 20451 14427 20457
rect 14369 20417 14381 20451
rect 14415 20417 14427 20451
rect 14369 20411 14427 20417
rect 15197 20451 15255 20457
rect 15197 20417 15209 20451
rect 15243 20448 15255 20451
rect 17126 20448 17132 20460
rect 15243 20420 17132 20448
rect 15243 20417 15255 20420
rect 15197 20411 15255 20417
rect 17126 20408 17132 20420
rect 17184 20408 17190 20460
rect 18046 20448 18052 20460
rect 18007 20420 18052 20448
rect 18046 20408 18052 20420
rect 18104 20408 18110 20460
rect 18233 20451 18291 20457
rect 18233 20417 18245 20451
rect 18279 20448 18291 20451
rect 18984 20448 19012 20476
rect 18279 20420 19012 20448
rect 19981 20451 20039 20457
rect 18279 20417 18291 20420
rect 18233 20411 18291 20417
rect 19981 20417 19993 20451
rect 20027 20448 20039 20451
rect 20088 20448 20116 20476
rect 20027 20420 20116 20448
rect 20257 20451 20315 20457
rect 20027 20417 20039 20420
rect 19981 20411 20039 20417
rect 20257 20417 20269 20451
rect 20303 20448 20315 20451
rect 20806 20448 20812 20460
rect 20303 20420 20812 20448
rect 20303 20417 20315 20420
rect 20257 20411 20315 20417
rect 15473 20383 15531 20389
rect 15473 20380 15485 20383
rect 14108 20352 15485 20380
rect 15473 20349 15485 20352
rect 15519 20380 15531 20383
rect 15654 20380 15660 20392
rect 15519 20352 15660 20380
rect 15519 20349 15531 20352
rect 15473 20343 15531 20349
rect 15654 20340 15660 20352
rect 15712 20340 15718 20392
rect 16390 20340 16396 20392
rect 16448 20380 16454 20392
rect 17497 20383 17555 20389
rect 17497 20380 17509 20383
rect 16448 20352 17509 20380
rect 16448 20340 16454 20352
rect 17497 20349 17509 20352
rect 17543 20380 17555 20383
rect 17770 20380 17776 20392
rect 17543 20352 17776 20380
rect 17543 20349 17555 20352
rect 17497 20343 17555 20349
rect 17770 20340 17776 20352
rect 17828 20340 17834 20392
rect 14093 20315 14151 20321
rect 14093 20312 14105 20315
rect 13832 20284 14105 20312
rect 13541 20275 13599 20281
rect 14093 20281 14105 20284
rect 14139 20281 14151 20315
rect 14093 20275 14151 20281
rect 16574 20272 16580 20324
rect 16632 20312 16638 20324
rect 18248 20312 18276 20411
rect 20806 20408 20812 20420
rect 20864 20408 20870 20460
rect 21100 20448 21128 20488
rect 21174 20476 21180 20528
rect 21232 20516 21238 20528
rect 22186 20516 22192 20528
rect 21232 20488 22192 20516
rect 21232 20476 21238 20488
rect 22186 20476 22192 20488
rect 22244 20476 22250 20528
rect 23658 20476 23664 20528
rect 23716 20516 23722 20528
rect 24946 20516 24952 20528
rect 23716 20488 24440 20516
rect 24907 20488 24952 20516
rect 23716 20476 23722 20488
rect 22002 20448 22008 20460
rect 21100 20420 22008 20448
rect 22002 20408 22008 20420
rect 22060 20408 22066 20460
rect 22094 20408 22100 20460
rect 22152 20448 22158 20460
rect 22278 20448 22284 20460
rect 22152 20420 22197 20448
rect 22239 20420 22284 20448
rect 22152 20408 22158 20420
rect 22278 20408 22284 20420
rect 22336 20408 22342 20460
rect 22462 20448 22468 20460
rect 22423 20420 22468 20448
rect 22462 20408 22468 20420
rect 22520 20408 22526 20460
rect 23014 20408 23020 20460
rect 23072 20448 23078 20460
rect 23109 20451 23167 20457
rect 23109 20448 23121 20451
rect 23072 20420 23121 20448
rect 23072 20408 23078 20420
rect 23109 20417 23121 20420
rect 23155 20417 23167 20451
rect 23934 20448 23940 20460
rect 23895 20420 23940 20448
rect 23109 20411 23167 20417
rect 23934 20408 23940 20420
rect 23992 20408 23998 20460
rect 24210 20448 24216 20460
rect 24171 20420 24216 20448
rect 24210 20408 24216 20420
rect 24268 20408 24274 20460
rect 24412 20457 24440 20488
rect 24946 20476 24952 20488
rect 25004 20476 25010 20528
rect 24397 20451 24455 20457
rect 24397 20417 24409 20451
rect 24443 20448 24455 20451
rect 25038 20448 25044 20460
rect 24443 20420 25044 20448
rect 24443 20417 24455 20420
rect 24397 20411 24455 20417
rect 25038 20408 25044 20420
rect 25096 20408 25102 20460
rect 25608 20448 25636 20556
rect 25774 20544 25780 20596
rect 25832 20584 25838 20596
rect 25885 20587 25943 20593
rect 25885 20584 25897 20587
rect 25832 20556 25897 20584
rect 25832 20544 25838 20556
rect 25885 20553 25897 20556
rect 25931 20553 25943 20587
rect 25885 20547 25943 20553
rect 29914 20544 29920 20596
rect 29972 20584 29978 20596
rect 30193 20587 30251 20593
rect 30193 20584 30205 20587
rect 29972 20556 30205 20584
rect 29972 20544 29978 20556
rect 30193 20553 30205 20556
rect 30239 20584 30251 20587
rect 30926 20584 30932 20596
rect 30239 20556 30932 20584
rect 30239 20553 30251 20556
rect 30193 20547 30251 20553
rect 30926 20544 30932 20556
rect 30984 20544 30990 20596
rect 33137 20587 33195 20593
rect 33137 20584 33149 20587
rect 31726 20556 33149 20584
rect 25685 20519 25743 20525
rect 25685 20485 25697 20519
rect 25731 20516 25743 20519
rect 26510 20516 26516 20528
rect 25731 20488 26516 20516
rect 25731 20485 25743 20488
rect 25685 20479 25743 20485
rect 26510 20476 26516 20488
rect 26568 20476 26574 20528
rect 26786 20476 26792 20528
rect 26844 20516 26850 20528
rect 27341 20519 27399 20525
rect 26844 20488 27200 20516
rect 26844 20476 26850 20488
rect 26694 20448 26700 20460
rect 25608 20420 26700 20448
rect 26694 20408 26700 20420
rect 26752 20448 26758 20460
rect 26878 20448 26884 20460
rect 26752 20420 26884 20448
rect 26752 20408 26758 20420
rect 26878 20408 26884 20420
rect 26936 20408 26942 20460
rect 27062 20448 27068 20460
rect 27023 20420 27068 20448
rect 27062 20408 27068 20420
rect 27120 20408 27126 20460
rect 27172 20457 27200 20488
rect 27341 20485 27353 20519
rect 27387 20516 27399 20519
rect 27706 20516 27712 20528
rect 27387 20488 27712 20516
rect 27387 20485 27399 20488
rect 27341 20479 27399 20485
rect 27706 20476 27712 20488
rect 27764 20476 27770 20528
rect 27982 20476 27988 20528
rect 28040 20516 28046 20528
rect 28040 20488 29132 20516
rect 28040 20476 28046 20488
rect 27158 20451 27216 20457
rect 27158 20417 27170 20451
rect 27204 20417 27216 20451
rect 27158 20411 27216 20417
rect 27433 20451 27491 20457
rect 27433 20417 27445 20451
rect 27479 20417 27491 20451
rect 27433 20411 27491 20417
rect 27571 20451 27629 20457
rect 27571 20417 27583 20451
rect 27617 20448 27629 20451
rect 28626 20448 28632 20460
rect 27617 20420 28632 20448
rect 27617 20417 27629 20420
rect 27571 20411 27629 20417
rect 22830 20380 22836 20392
rect 22066 20352 22836 20380
rect 16632 20284 18276 20312
rect 19076 20284 19380 20312
rect 16632 20272 16638 20284
rect 9122 20244 9128 20256
rect 8956 20216 9128 20244
rect 9122 20204 9128 20216
rect 9180 20244 9186 20256
rect 15838 20244 15844 20256
rect 9180 20216 15844 20244
rect 9180 20204 9186 20216
rect 15838 20204 15844 20216
rect 15896 20204 15902 20256
rect 16850 20244 16856 20256
rect 16811 20216 16856 20244
rect 16850 20204 16856 20216
rect 16908 20204 16914 20256
rect 19076 20253 19104 20284
rect 19061 20247 19119 20253
rect 19061 20213 19073 20247
rect 19107 20213 19119 20247
rect 19352 20244 19380 20284
rect 20622 20272 20628 20324
rect 20680 20312 20686 20324
rect 22066 20312 22094 20352
rect 22830 20340 22836 20352
rect 22888 20340 22894 20392
rect 23290 20340 23296 20392
rect 23348 20380 23354 20392
rect 23348 20352 23796 20380
rect 23348 20340 23354 20352
rect 20680 20284 22094 20312
rect 22189 20315 22247 20321
rect 20680 20272 20686 20284
rect 22189 20281 22201 20315
rect 22235 20312 22247 20315
rect 23474 20312 23480 20324
rect 22235 20284 23480 20312
rect 22235 20281 22247 20284
rect 22189 20275 22247 20281
rect 23474 20272 23480 20284
rect 23532 20272 23538 20324
rect 23768 20312 23796 20352
rect 24029 20315 24087 20321
rect 24029 20312 24041 20315
rect 23768 20284 24041 20312
rect 24029 20281 24041 20284
rect 24075 20281 24087 20315
rect 24029 20275 24087 20281
rect 24121 20315 24179 20321
rect 24121 20281 24133 20315
rect 24167 20312 24179 20315
rect 25590 20312 25596 20324
rect 24167 20284 25596 20312
rect 24167 20281 24179 20284
rect 24121 20275 24179 20281
rect 25590 20272 25596 20284
rect 25648 20272 25654 20324
rect 26326 20312 26332 20324
rect 25884 20284 26332 20312
rect 20993 20247 21051 20253
rect 20993 20244 21005 20247
rect 19352 20216 21005 20244
rect 19061 20207 19119 20213
rect 20993 20213 21005 20216
rect 21039 20213 21051 20247
rect 20993 20207 21051 20213
rect 22370 20204 22376 20256
rect 22428 20244 22434 20256
rect 23753 20247 23811 20253
rect 23753 20244 23765 20247
rect 22428 20216 23765 20244
rect 22428 20204 22434 20216
rect 23753 20213 23765 20216
rect 23799 20213 23811 20247
rect 23753 20207 23811 20213
rect 25041 20247 25099 20253
rect 25041 20213 25053 20247
rect 25087 20244 25099 20247
rect 25498 20244 25504 20256
rect 25087 20216 25504 20244
rect 25087 20213 25099 20216
rect 25041 20207 25099 20213
rect 25498 20204 25504 20216
rect 25556 20204 25562 20256
rect 25884 20253 25912 20284
rect 26326 20272 26332 20284
rect 26384 20272 26390 20324
rect 27448 20312 27476 20411
rect 28626 20408 28632 20420
rect 28684 20408 28690 20460
rect 28994 20448 29000 20460
rect 28955 20420 29000 20448
rect 28994 20408 29000 20420
rect 29052 20408 29058 20460
rect 29104 20448 29132 20488
rect 29178 20476 29184 20528
rect 29236 20516 29242 20528
rect 30098 20516 30104 20528
rect 29236 20488 30104 20516
rect 29236 20476 29242 20488
rect 30098 20476 30104 20488
rect 30156 20516 30162 20528
rect 31726 20516 31754 20556
rect 33137 20553 33149 20556
rect 33183 20553 33195 20587
rect 33137 20547 33195 20553
rect 35434 20544 35440 20596
rect 35492 20584 35498 20596
rect 35529 20587 35587 20593
rect 35529 20584 35541 20587
rect 35492 20556 35541 20584
rect 35492 20544 35498 20556
rect 35529 20553 35541 20556
rect 35575 20553 35587 20587
rect 35529 20547 35587 20553
rect 30156 20488 31754 20516
rect 32677 20519 32735 20525
rect 30156 20476 30162 20488
rect 32677 20485 32689 20519
rect 32723 20516 32735 20519
rect 33226 20516 33232 20528
rect 32723 20488 33232 20516
rect 32723 20485 32735 20488
rect 32677 20479 32735 20485
rect 33226 20476 33232 20488
rect 33284 20476 33290 20528
rect 33870 20516 33876 20528
rect 33520 20488 33876 20516
rect 31205 20451 31263 20457
rect 31205 20448 31217 20451
rect 29104 20420 31217 20448
rect 31205 20417 31217 20420
rect 31251 20417 31263 20451
rect 31205 20411 31263 20417
rect 31389 20451 31447 20457
rect 31389 20417 31401 20451
rect 31435 20448 31447 20451
rect 32030 20448 32036 20460
rect 31435 20420 32036 20448
rect 31435 20417 31447 20420
rect 31389 20411 31447 20417
rect 28074 20340 28080 20392
rect 28132 20380 28138 20392
rect 28718 20380 28724 20392
rect 28132 20352 28724 20380
rect 28132 20340 28138 20352
rect 28718 20340 28724 20352
rect 28776 20340 28782 20392
rect 31220 20380 31248 20411
rect 32030 20408 32036 20420
rect 32088 20408 32094 20460
rect 32122 20408 32128 20460
rect 32180 20448 32186 20460
rect 32220 20451 32278 20457
rect 32220 20448 32232 20451
rect 32180 20420 32232 20448
rect 32180 20408 32186 20420
rect 32220 20417 32232 20420
rect 32266 20448 32278 20451
rect 32490 20448 32496 20460
rect 32266 20420 32353 20448
rect 32451 20420 32496 20448
rect 32266 20417 32278 20420
rect 32220 20411 32278 20417
rect 31662 20380 31668 20392
rect 31220 20352 31668 20380
rect 31662 20340 31668 20352
rect 31720 20340 31726 20392
rect 32325 20380 32353 20420
rect 32490 20408 32496 20420
rect 32548 20408 32554 20460
rect 33520 20457 33548 20488
rect 33870 20476 33876 20488
rect 33928 20516 33934 20528
rect 33928 20488 34468 20516
rect 33928 20476 33934 20488
rect 34440 20457 34468 20488
rect 34790 20476 34796 20528
rect 34848 20516 34854 20528
rect 34977 20519 35035 20525
rect 34977 20516 34989 20519
rect 34848 20488 34989 20516
rect 34848 20476 34854 20488
rect 34977 20485 34989 20488
rect 35023 20485 35035 20519
rect 36357 20519 36415 20525
rect 36357 20516 36369 20519
rect 34977 20479 35035 20485
rect 35728 20488 36369 20516
rect 33505 20451 33563 20457
rect 33505 20417 33517 20451
rect 33551 20417 33563 20451
rect 33505 20411 33563 20417
rect 34241 20451 34299 20457
rect 34241 20417 34253 20451
rect 34287 20417 34299 20451
rect 34241 20411 34299 20417
rect 34425 20451 34483 20457
rect 34425 20417 34437 20451
rect 34471 20417 34483 20451
rect 34425 20411 34483 20417
rect 33318 20380 33324 20392
rect 32325 20352 33324 20380
rect 33318 20340 33324 20352
rect 33376 20340 33382 20392
rect 33597 20383 33655 20389
rect 33597 20349 33609 20383
rect 33643 20380 33655 20383
rect 34256 20380 34284 20411
rect 34698 20408 34704 20460
rect 34756 20448 34762 20460
rect 35728 20457 35756 20488
rect 36357 20485 36369 20488
rect 36403 20485 36415 20519
rect 36357 20479 36415 20485
rect 35713 20451 35771 20457
rect 35713 20448 35725 20451
rect 34756 20420 35725 20448
rect 34756 20408 34762 20420
rect 35713 20417 35725 20420
rect 35759 20417 35771 20451
rect 36170 20448 36176 20460
rect 36131 20420 36176 20448
rect 35713 20411 35771 20417
rect 36170 20408 36176 20420
rect 36228 20408 36234 20460
rect 33643 20352 35112 20380
rect 33643 20349 33655 20352
rect 33597 20343 33655 20349
rect 29178 20312 29184 20324
rect 27448 20284 29184 20312
rect 29178 20272 29184 20284
rect 29236 20272 29242 20324
rect 34977 20315 35035 20321
rect 34977 20312 34989 20315
rect 32600 20284 34989 20312
rect 32600 20256 32628 20284
rect 34977 20281 34989 20284
rect 35023 20281 35035 20315
rect 35084 20312 35112 20352
rect 35342 20340 35348 20392
rect 35400 20380 35406 20392
rect 35437 20383 35495 20389
rect 35437 20380 35449 20383
rect 35400 20352 35449 20380
rect 35400 20340 35406 20352
rect 35437 20349 35449 20352
rect 35483 20380 35495 20383
rect 35986 20380 35992 20392
rect 35483 20352 35992 20380
rect 35483 20349 35495 20352
rect 35437 20343 35495 20349
rect 35986 20340 35992 20352
rect 36044 20340 36050 20392
rect 36541 20315 36599 20321
rect 36541 20312 36553 20315
rect 35084 20284 36553 20312
rect 34977 20275 35035 20281
rect 36541 20281 36553 20284
rect 36587 20281 36599 20315
rect 36541 20275 36599 20281
rect 25869 20247 25927 20253
rect 25869 20213 25881 20247
rect 25915 20213 25927 20247
rect 26050 20244 26056 20256
rect 26011 20216 26056 20244
rect 25869 20207 25927 20213
rect 26050 20204 26056 20216
rect 26108 20204 26114 20256
rect 27706 20204 27712 20256
rect 27764 20244 27770 20256
rect 31573 20247 31631 20253
rect 27764 20216 27809 20244
rect 27764 20204 27770 20216
rect 31573 20213 31585 20247
rect 31619 20244 31631 20247
rect 31754 20244 31760 20256
rect 31619 20216 31760 20244
rect 31619 20213 31631 20216
rect 31573 20207 31631 20213
rect 31754 20204 31760 20216
rect 31812 20204 31818 20256
rect 32582 20244 32588 20256
rect 32543 20216 32588 20244
rect 32582 20204 32588 20216
rect 32640 20204 32646 20256
rect 32766 20204 32772 20256
rect 32824 20244 32830 20256
rect 33781 20247 33839 20253
rect 33781 20244 33793 20247
rect 32824 20216 33793 20244
rect 32824 20204 32830 20216
rect 33781 20213 33793 20216
rect 33827 20213 33839 20247
rect 34238 20244 34244 20256
rect 34151 20216 34244 20244
rect 33781 20207 33839 20213
rect 34238 20204 34244 20216
rect 34296 20244 34302 20256
rect 35526 20244 35532 20256
rect 34296 20216 35532 20244
rect 34296 20204 34302 20216
rect 35526 20204 35532 20216
rect 35584 20204 35590 20256
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 7742 20040 7748 20052
rect 7703 20012 7748 20040
rect 7742 20000 7748 20012
rect 7800 20000 7806 20052
rect 7926 20000 7932 20052
rect 7984 20040 7990 20052
rect 19429 20043 19487 20049
rect 7984 20012 13676 20040
rect 7984 20000 7990 20012
rect 9122 19972 9128 19984
rect 8036 19944 9128 19972
rect 7926 19904 7932 19916
rect 7887 19876 7932 19904
rect 7926 19864 7932 19876
rect 7984 19864 7990 19916
rect 8036 19913 8064 19944
rect 9122 19932 9128 19944
rect 9180 19932 9186 19984
rect 10042 19972 10048 19984
rect 9508 19944 10048 19972
rect 8021 19907 8079 19913
rect 8021 19873 8033 19907
rect 8067 19873 8079 19907
rect 8386 19904 8392 19916
rect 8347 19876 8392 19904
rect 8021 19867 8079 19873
rect 8386 19864 8392 19876
rect 8444 19864 8450 19916
rect 9508 19913 9536 19944
rect 10042 19932 10048 19944
rect 10100 19972 10106 19984
rect 10962 19972 10968 19984
rect 10100 19944 10968 19972
rect 10100 19932 10106 19944
rect 10962 19932 10968 19944
rect 11020 19932 11026 19984
rect 13446 19972 13452 19984
rect 12452 19944 13452 19972
rect 9493 19907 9551 19913
rect 9493 19873 9505 19907
rect 9539 19873 9551 19907
rect 11974 19904 11980 19916
rect 9493 19867 9551 19873
rect 10888 19876 11980 19904
rect 8297 19839 8355 19845
rect 8297 19805 8309 19839
rect 8343 19836 8355 19839
rect 8754 19836 8760 19848
rect 8343 19808 8760 19836
rect 8343 19805 8355 19808
rect 8297 19799 8355 19805
rect 8754 19796 8760 19808
rect 8812 19796 8818 19848
rect 10888 19845 10916 19876
rect 11974 19864 11980 19876
rect 12032 19864 12038 19916
rect 12342 19904 12348 19916
rect 12303 19876 12348 19904
rect 12342 19864 12348 19876
rect 12400 19864 12406 19916
rect 12452 19913 12480 19944
rect 13446 19932 13452 19944
rect 13504 19932 13510 19984
rect 12437 19907 12495 19913
rect 12437 19873 12449 19907
rect 12483 19873 12495 19907
rect 12618 19904 12624 19916
rect 12579 19876 12624 19904
rect 12437 19867 12495 19873
rect 12618 19864 12624 19876
rect 12676 19864 12682 19916
rect 13648 19904 13676 20012
rect 19429 20009 19441 20043
rect 19475 20040 19487 20043
rect 20070 20040 20076 20052
rect 19475 20012 20076 20040
rect 19475 20009 19487 20012
rect 19429 20003 19487 20009
rect 20070 20000 20076 20012
rect 20128 20000 20134 20052
rect 20533 20043 20591 20049
rect 20533 20009 20545 20043
rect 20579 20040 20591 20043
rect 22094 20040 22100 20052
rect 20579 20012 22100 20040
rect 20579 20009 20591 20012
rect 20533 20003 20591 20009
rect 22094 20000 22100 20012
rect 22152 20000 22158 20052
rect 23658 20040 23664 20052
rect 23619 20012 23664 20040
rect 23658 20000 23664 20012
rect 23716 20000 23722 20052
rect 23753 20043 23811 20049
rect 23753 20009 23765 20043
rect 23799 20040 23811 20043
rect 24210 20040 24216 20052
rect 23799 20012 24216 20040
rect 23799 20009 23811 20012
rect 23753 20003 23811 20009
rect 24210 20000 24216 20012
rect 24268 20000 24274 20052
rect 24762 20000 24768 20052
rect 24820 20040 24826 20052
rect 28261 20043 28319 20049
rect 24820 20012 27016 20040
rect 24820 20000 24826 20012
rect 15749 19975 15807 19981
rect 15749 19941 15761 19975
rect 15795 19941 15807 19975
rect 15749 19935 15807 19941
rect 15764 19904 15792 19935
rect 17494 19932 17500 19984
rect 17552 19972 17558 19984
rect 17552 19944 20760 19972
rect 17552 19932 17558 19944
rect 16114 19904 16120 19916
rect 13372 19876 14504 19904
rect 15764 19876 16120 19904
rect 9217 19839 9275 19845
rect 9217 19805 9229 19839
rect 9263 19805 9275 19839
rect 9217 19799 9275 19805
rect 10781 19839 10839 19845
rect 10781 19805 10793 19839
rect 10827 19805 10839 19839
rect 10781 19799 10839 19805
rect 10873 19839 10931 19845
rect 10873 19805 10885 19839
rect 10919 19805 10931 19839
rect 10873 19799 10931 19805
rect 10965 19836 11023 19842
rect 10965 19802 10977 19836
rect 11011 19802 11023 19836
rect 9232 19768 9260 19799
rect 10410 19768 10416 19780
rect 8220 19740 10416 19768
rect 8220 19709 8248 19740
rect 10410 19728 10416 19740
rect 10468 19728 10474 19780
rect 10796 19768 10824 19799
rect 10965 19796 11023 19802
rect 11125 19839 11183 19845
rect 11125 19805 11137 19839
rect 11171 19836 11183 19839
rect 11330 19836 11336 19848
rect 11171 19830 11192 19836
rect 11256 19830 11336 19836
rect 11171 19808 11336 19830
rect 11171 19805 11284 19808
rect 11125 19802 11284 19805
rect 11125 19799 11183 19802
rect 11330 19796 11336 19808
rect 11388 19796 11394 19848
rect 12529 19839 12587 19845
rect 12529 19805 12541 19839
rect 12575 19836 12587 19839
rect 12802 19836 12808 19848
rect 12575 19808 12808 19836
rect 12575 19805 12587 19808
rect 12529 19799 12587 19805
rect 12802 19796 12808 19808
rect 12860 19796 12866 19848
rect 13372 19845 13400 19876
rect 13357 19839 13415 19845
rect 13357 19805 13369 19839
rect 13403 19805 13415 19839
rect 14366 19836 14372 19848
rect 14327 19808 14372 19836
rect 13357 19799 13415 19805
rect 14366 19796 14372 19808
rect 14424 19796 14430 19848
rect 14476 19836 14504 19876
rect 16114 19864 16120 19876
rect 16172 19904 16178 19916
rect 16209 19907 16267 19913
rect 16209 19904 16221 19907
rect 16172 19876 16221 19904
rect 16172 19864 16178 19876
rect 16209 19873 16221 19876
rect 16255 19873 16267 19907
rect 16482 19904 16488 19916
rect 16443 19876 16488 19904
rect 16209 19867 16267 19873
rect 16482 19864 16488 19876
rect 16540 19864 16546 19916
rect 17862 19904 17868 19916
rect 17823 19876 17868 19904
rect 17862 19864 17868 19876
rect 17920 19864 17926 19916
rect 18141 19907 18199 19913
rect 18141 19873 18153 19907
rect 18187 19904 18199 19907
rect 18230 19904 18236 19916
rect 18187 19876 18236 19904
rect 18187 19873 18199 19876
rect 18141 19867 18199 19873
rect 18230 19864 18236 19876
rect 18288 19904 18294 19916
rect 18288 19876 20392 19904
rect 18288 19864 18294 19876
rect 15838 19836 15844 19848
rect 14476 19808 15844 19836
rect 15838 19796 15844 19808
rect 15896 19796 15902 19848
rect 17954 19796 17960 19848
rect 18012 19836 18018 19848
rect 19978 19836 19984 19848
rect 18012 19808 19840 19836
rect 19939 19808 19984 19836
rect 18012 19796 18018 19808
rect 10704 19740 10824 19768
rect 8205 19703 8263 19709
rect 8205 19669 8217 19703
rect 8251 19669 8263 19703
rect 10502 19700 10508 19712
rect 10463 19672 10508 19700
rect 8205 19663 8263 19669
rect 10502 19660 10508 19672
rect 10560 19660 10566 19712
rect 10594 19660 10600 19712
rect 10652 19700 10658 19712
rect 10704 19700 10732 19740
rect 10652 19672 10732 19700
rect 10980 19700 11008 19796
rect 14274 19728 14280 19780
rect 14332 19768 14338 19780
rect 14614 19771 14672 19777
rect 14614 19768 14626 19771
rect 14332 19740 14626 19768
rect 14332 19728 14338 19740
rect 14614 19737 14626 19740
rect 14660 19737 14672 19771
rect 19334 19768 19340 19780
rect 19295 19740 19340 19768
rect 14614 19731 14672 19737
rect 19334 19728 19340 19740
rect 19392 19728 19398 19780
rect 19812 19768 19840 19808
rect 19978 19796 19984 19808
rect 20036 19796 20042 19848
rect 20364 19845 20392 19876
rect 20349 19839 20407 19845
rect 20349 19805 20361 19839
rect 20395 19836 20407 19839
rect 20622 19836 20628 19848
rect 20395 19808 20628 19836
rect 20395 19805 20407 19808
rect 20349 19799 20407 19805
rect 20622 19796 20628 19808
rect 20680 19796 20686 19848
rect 20732 19836 20760 19944
rect 26142 19932 26148 19984
rect 26200 19972 26206 19984
rect 26878 19972 26884 19984
rect 26200 19944 26740 19972
rect 26839 19944 26884 19972
rect 26200 19932 26206 19944
rect 20990 19904 20996 19916
rect 20951 19876 20996 19904
rect 20990 19864 20996 19876
rect 21048 19864 21054 19916
rect 22186 19864 22192 19916
rect 22244 19904 22250 19916
rect 23842 19904 23848 19916
rect 22244 19876 22508 19904
rect 23803 19876 23848 19904
rect 22244 19864 22250 19876
rect 21174 19836 21180 19848
rect 20732 19808 21180 19836
rect 21174 19796 21180 19808
rect 21232 19796 21238 19848
rect 21269 19839 21327 19845
rect 21269 19805 21281 19839
rect 21315 19836 21327 19839
rect 22370 19836 22376 19848
rect 21315 19808 22376 19836
rect 21315 19805 21327 19808
rect 21269 19799 21327 19805
rect 22370 19796 22376 19808
rect 22428 19796 22434 19848
rect 22480 19845 22508 19876
rect 23842 19864 23848 19876
rect 23900 19864 23906 19916
rect 24762 19904 24768 19916
rect 24723 19876 24768 19904
rect 24762 19864 24768 19876
rect 24820 19864 24826 19916
rect 25774 19864 25780 19916
rect 25832 19904 25838 19916
rect 26712 19904 26740 19944
rect 26878 19932 26884 19944
rect 26936 19932 26942 19984
rect 26988 19972 27016 20012
rect 28261 20009 28273 20043
rect 28307 20040 28319 20043
rect 28350 20040 28356 20052
rect 28307 20012 28356 20040
rect 28307 20009 28319 20012
rect 28261 20003 28319 20009
rect 28350 20000 28356 20012
rect 28408 20000 28414 20052
rect 28718 20000 28724 20052
rect 28776 20040 28782 20052
rect 29549 20043 29607 20049
rect 29549 20040 29561 20043
rect 28776 20012 29561 20040
rect 28776 20000 28782 20012
rect 29549 20009 29561 20012
rect 29595 20009 29607 20043
rect 29549 20003 29607 20009
rect 31481 20043 31539 20049
rect 31481 20009 31493 20043
rect 31527 20040 31539 20043
rect 32122 20040 32128 20052
rect 31527 20012 32128 20040
rect 31527 20009 31539 20012
rect 31481 20003 31539 20009
rect 32122 20000 32128 20012
rect 32180 20000 32186 20052
rect 32766 20040 32772 20052
rect 32727 20012 32772 20040
rect 32766 20000 32772 20012
rect 32824 20000 32830 20052
rect 34885 20043 34943 20049
rect 34885 20009 34897 20043
rect 34931 20040 34943 20043
rect 36170 20040 36176 20052
rect 34931 20012 36176 20040
rect 34931 20009 34943 20012
rect 34885 20003 34943 20009
rect 36170 20000 36176 20012
rect 36228 20000 36234 20052
rect 29270 19972 29276 19984
rect 26988 19944 29276 19972
rect 29270 19932 29276 19944
rect 29328 19932 29334 19984
rect 29380 19944 32628 19972
rect 29380 19904 29408 19944
rect 32030 19904 32036 19916
rect 25832 19876 26280 19904
rect 26712 19876 29408 19904
rect 31496 19876 32036 19904
rect 25832 19864 25838 19876
rect 22465 19839 22523 19845
rect 22465 19805 22477 19839
rect 22511 19805 22523 19839
rect 22830 19836 22836 19848
rect 22743 19808 22836 19836
rect 22465 19799 22523 19805
rect 22830 19796 22836 19808
rect 22888 19836 22894 19848
rect 23382 19836 23388 19848
rect 22888 19808 23388 19836
rect 22888 19796 22894 19808
rect 23382 19796 23388 19808
rect 23440 19796 23446 19848
rect 23566 19836 23572 19848
rect 23527 19808 23572 19836
rect 23566 19796 23572 19808
rect 23624 19796 23630 19848
rect 23934 19796 23940 19848
rect 23992 19836 23998 19848
rect 24486 19836 24492 19848
rect 23992 19808 24492 19836
rect 23992 19796 23998 19808
rect 24486 19796 24492 19808
rect 24544 19836 24550 19848
rect 24581 19839 24639 19845
rect 24581 19836 24593 19839
rect 24544 19808 24593 19836
rect 24544 19796 24550 19808
rect 24581 19805 24593 19808
rect 24627 19805 24639 19839
rect 24581 19799 24639 19805
rect 24673 19839 24731 19845
rect 24673 19805 24685 19839
rect 24719 19805 24731 19839
rect 24673 19799 24731 19805
rect 20162 19768 20168 19780
rect 19812 19740 20168 19768
rect 20162 19728 20168 19740
rect 20220 19728 20226 19780
rect 20257 19771 20315 19777
rect 20257 19737 20269 19771
rect 20303 19768 20315 19771
rect 22646 19768 22652 19780
rect 20303 19740 22048 19768
rect 22607 19740 22652 19768
rect 20303 19737 20315 19740
rect 20257 19731 20315 19737
rect 11054 19700 11060 19712
rect 10980 19672 11060 19700
rect 10652 19660 10658 19672
rect 11054 19660 11060 19672
rect 11112 19660 11118 19712
rect 12161 19703 12219 19709
rect 12161 19669 12173 19703
rect 12207 19700 12219 19703
rect 12618 19700 12624 19712
rect 12207 19672 12624 19700
rect 12207 19669 12219 19672
rect 12161 19663 12219 19669
rect 12618 19660 12624 19672
rect 12676 19660 12682 19712
rect 13446 19700 13452 19712
rect 13359 19672 13452 19700
rect 13446 19660 13452 19672
rect 13504 19700 13510 19712
rect 15654 19700 15660 19712
rect 13504 19672 15660 19700
rect 13504 19660 13510 19672
rect 15654 19660 15660 19672
rect 15712 19700 15718 19712
rect 20530 19700 20536 19712
rect 15712 19672 20536 19700
rect 15712 19660 15718 19672
rect 20530 19660 20536 19672
rect 20588 19660 20594 19712
rect 22020 19709 22048 19740
rect 22646 19728 22652 19740
rect 22704 19728 22710 19780
rect 22738 19728 22744 19780
rect 22796 19768 22802 19780
rect 22796 19740 22841 19768
rect 22796 19728 22802 19740
rect 22922 19728 22928 19780
rect 22980 19768 22986 19780
rect 24688 19768 24716 19799
rect 24854 19796 24860 19848
rect 24912 19836 24918 19848
rect 24912 19808 24957 19836
rect 24912 19796 24918 19808
rect 25038 19796 25044 19848
rect 25096 19836 25102 19848
rect 25096 19808 25141 19836
rect 25096 19796 25102 19808
rect 25958 19796 25964 19848
rect 26016 19836 26022 19848
rect 26252 19845 26280 19876
rect 26053 19839 26111 19845
rect 26053 19836 26065 19839
rect 26016 19808 26065 19836
rect 26016 19796 26022 19808
rect 26053 19805 26065 19808
rect 26099 19805 26111 19839
rect 26053 19799 26111 19805
rect 26237 19839 26295 19845
rect 26237 19805 26249 19839
rect 26283 19805 26295 19839
rect 26237 19799 26295 19805
rect 22980 19740 24716 19768
rect 26252 19768 26280 19799
rect 26326 19796 26332 19848
rect 26384 19836 26390 19848
rect 27157 19839 27215 19845
rect 27157 19836 27169 19839
rect 26384 19808 27169 19836
rect 26384 19796 26390 19808
rect 27157 19805 27169 19808
rect 27203 19805 27215 19839
rect 28442 19836 28448 19848
rect 27157 19799 27215 19805
rect 28092 19808 28448 19836
rect 28092 19777 28120 19808
rect 28442 19796 28448 19808
rect 28500 19796 28506 19848
rect 28994 19836 29000 19848
rect 28828 19808 29000 19836
rect 26881 19771 26939 19777
rect 26881 19768 26893 19771
rect 26252 19740 26893 19768
rect 22980 19728 22986 19740
rect 26881 19737 26893 19740
rect 26927 19737 26939 19771
rect 26881 19731 26939 19737
rect 28077 19771 28135 19777
rect 28077 19737 28089 19771
rect 28123 19737 28135 19771
rect 28077 19731 28135 19737
rect 28293 19771 28351 19777
rect 28293 19737 28305 19771
rect 28339 19768 28351 19771
rect 28828 19768 28856 19808
rect 28994 19796 29000 19808
rect 29052 19796 29058 19848
rect 29362 19796 29368 19848
rect 29420 19836 29426 19848
rect 29549 19839 29607 19845
rect 29549 19836 29561 19839
rect 29420 19808 29561 19836
rect 29420 19796 29426 19808
rect 29549 19805 29561 19808
rect 29595 19805 29607 19839
rect 29730 19836 29736 19848
rect 29691 19808 29736 19836
rect 29549 19799 29607 19805
rect 29730 19796 29736 19808
rect 29788 19796 29794 19848
rect 30558 19836 30564 19848
rect 30519 19808 30564 19836
rect 30558 19796 30564 19808
rect 30616 19796 30622 19848
rect 30745 19839 30803 19845
rect 30745 19805 30757 19839
rect 30791 19836 30803 19839
rect 31110 19836 31116 19848
rect 30791 19808 31116 19836
rect 30791 19805 30803 19808
rect 30745 19799 30803 19805
rect 31110 19796 31116 19808
rect 31168 19796 31174 19848
rect 31496 19845 31524 19876
rect 32030 19864 32036 19876
rect 32088 19864 32094 19916
rect 31481 19839 31539 19845
rect 31481 19805 31493 19839
rect 31527 19805 31539 19839
rect 31662 19836 31668 19848
rect 31623 19808 31668 19836
rect 31481 19799 31539 19805
rect 31662 19796 31668 19808
rect 31720 19796 31726 19848
rect 32600 19845 32628 19944
rect 34790 19932 34796 19984
rect 34848 19972 34854 19984
rect 35437 19975 35495 19981
rect 35437 19972 35449 19975
rect 34848 19944 35449 19972
rect 34848 19932 34854 19944
rect 35437 19941 35449 19944
rect 35483 19941 35495 19975
rect 35437 19935 35495 19941
rect 32861 19907 32919 19913
rect 32861 19873 32873 19907
rect 32907 19904 32919 19907
rect 34238 19904 34244 19916
rect 32907 19876 34244 19904
rect 32907 19873 32919 19876
rect 32861 19867 32919 19873
rect 34238 19864 34244 19876
rect 34296 19864 34302 19916
rect 35250 19864 35256 19916
rect 35308 19904 35314 19916
rect 35529 19907 35587 19913
rect 35529 19904 35541 19907
rect 35308 19876 35541 19904
rect 35308 19864 35314 19876
rect 35529 19873 35541 19876
rect 35575 19873 35587 19907
rect 35529 19867 35587 19873
rect 32585 19839 32643 19845
rect 32585 19805 32597 19839
rect 32631 19805 32643 19839
rect 32585 19799 32643 19805
rect 35066 19839 35124 19845
rect 35066 19805 35078 19839
rect 35112 19836 35124 19839
rect 35342 19836 35348 19848
rect 35112 19808 35348 19836
rect 35112 19805 35124 19808
rect 35066 19799 35124 19805
rect 35342 19796 35348 19808
rect 35400 19796 35406 19848
rect 28339 19740 28856 19768
rect 28339 19737 28351 19740
rect 28293 19731 28351 19737
rect 28902 19728 28908 19780
rect 28960 19768 28966 19780
rect 34330 19768 34336 19780
rect 28960 19740 34336 19768
rect 28960 19728 28966 19740
rect 34330 19728 34336 19740
rect 34388 19728 34394 19780
rect 22005 19703 22063 19709
rect 22005 19669 22017 19703
rect 22051 19669 22063 19703
rect 23014 19700 23020 19712
rect 22975 19672 23020 19700
rect 22005 19663 22063 19669
rect 23014 19660 23020 19672
rect 23072 19660 23078 19712
rect 23474 19660 23480 19712
rect 23532 19700 23538 19712
rect 24397 19703 24455 19709
rect 24397 19700 24409 19703
rect 23532 19672 24409 19700
rect 23532 19660 23538 19672
rect 24397 19669 24409 19672
rect 24443 19669 24455 19703
rect 24397 19663 24455 19669
rect 25774 19660 25780 19712
rect 25832 19700 25838 19712
rect 26421 19703 26479 19709
rect 26421 19700 26433 19703
rect 25832 19672 26433 19700
rect 25832 19660 25838 19672
rect 26421 19669 26433 19672
rect 26467 19669 26479 19703
rect 26421 19663 26479 19669
rect 26510 19660 26516 19712
rect 26568 19700 26574 19712
rect 27065 19703 27123 19709
rect 27065 19700 27077 19703
rect 26568 19672 27077 19700
rect 26568 19660 26574 19672
rect 27065 19669 27077 19672
rect 27111 19700 27123 19703
rect 28166 19700 28172 19712
rect 27111 19672 28172 19700
rect 27111 19669 27123 19672
rect 27065 19663 27123 19669
rect 28166 19660 28172 19672
rect 28224 19660 28230 19712
rect 28442 19700 28448 19712
rect 28403 19672 28448 19700
rect 28442 19660 28448 19672
rect 28500 19660 28506 19712
rect 29546 19660 29552 19712
rect 29604 19700 29610 19712
rect 30466 19700 30472 19712
rect 29604 19672 30472 19700
rect 29604 19660 29610 19672
rect 30466 19660 30472 19672
rect 30524 19660 30530 19712
rect 30745 19703 30803 19709
rect 30745 19669 30757 19703
rect 30791 19700 30803 19703
rect 31018 19700 31024 19712
rect 30791 19672 31024 19700
rect 30791 19669 30803 19672
rect 30745 19663 30803 19669
rect 31018 19660 31024 19672
rect 31076 19660 31082 19712
rect 32398 19700 32404 19712
rect 32359 19672 32404 19700
rect 32398 19660 32404 19672
rect 32456 19660 32462 19712
rect 33042 19660 33048 19712
rect 33100 19700 33106 19712
rect 34974 19700 34980 19712
rect 33100 19672 34980 19700
rect 33100 19660 33106 19672
rect 34974 19660 34980 19672
rect 35032 19660 35038 19712
rect 35069 19703 35127 19709
rect 35069 19669 35081 19703
rect 35115 19700 35127 19703
rect 35434 19700 35440 19712
rect 35115 19672 35440 19700
rect 35115 19669 35127 19672
rect 35069 19663 35127 19669
rect 35434 19660 35440 19672
rect 35492 19660 35498 19712
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 9122 19496 9128 19508
rect 9083 19468 9128 19496
rect 9122 19456 9128 19468
rect 9180 19456 9186 19508
rect 10137 19499 10195 19505
rect 10137 19465 10149 19499
rect 10183 19496 10195 19499
rect 10318 19496 10324 19508
rect 10183 19468 10324 19496
rect 10183 19465 10195 19468
rect 10137 19459 10195 19465
rect 10318 19456 10324 19468
rect 10376 19456 10382 19508
rect 14283 19499 14341 19505
rect 14283 19496 14295 19499
rect 10520 19468 14295 19496
rect 7282 19388 7288 19440
rect 7340 19428 7346 19440
rect 9398 19428 9404 19440
rect 7340 19400 9404 19428
rect 7340 19388 7346 19400
rect 7760 19369 7788 19400
rect 9398 19388 9404 19400
rect 9456 19388 9462 19440
rect 10226 19388 10232 19440
rect 10284 19428 10290 19440
rect 10520 19428 10548 19468
rect 14283 19465 14295 19468
rect 14329 19465 14341 19499
rect 14283 19459 14341 19465
rect 15473 19499 15531 19505
rect 15473 19465 15485 19499
rect 15519 19496 15531 19499
rect 15930 19496 15936 19508
rect 15519 19468 15936 19496
rect 15519 19465 15531 19468
rect 15473 19459 15531 19465
rect 15930 19456 15936 19468
rect 15988 19496 15994 19508
rect 16482 19496 16488 19508
rect 15988 19468 16488 19496
rect 15988 19456 15994 19468
rect 16482 19456 16488 19468
rect 16540 19456 16546 19508
rect 17126 19456 17132 19508
rect 17184 19496 17190 19508
rect 18325 19499 18383 19505
rect 18325 19496 18337 19499
rect 17184 19468 18337 19496
rect 17184 19456 17190 19468
rect 18325 19465 18337 19468
rect 18371 19465 18383 19499
rect 18325 19459 18383 19465
rect 19429 19499 19487 19505
rect 19429 19465 19441 19499
rect 19475 19496 19487 19499
rect 19978 19496 19984 19508
rect 19475 19468 19984 19496
rect 19475 19465 19487 19468
rect 19429 19459 19487 19465
rect 19978 19456 19984 19468
rect 20036 19456 20042 19508
rect 20346 19496 20352 19508
rect 20088 19468 20352 19496
rect 10284 19400 10548 19428
rect 10284 19388 10290 19400
rect 8018 19369 8024 19372
rect 7745 19363 7803 19369
rect 7745 19329 7757 19363
rect 7791 19329 7803 19363
rect 7745 19323 7803 19329
rect 8012 19323 8024 19369
rect 8076 19360 8082 19372
rect 10318 19360 10324 19372
rect 8076 19332 8112 19360
rect 10279 19332 10324 19360
rect 8018 19320 8024 19323
rect 8076 19320 8082 19332
rect 10318 19320 10324 19332
rect 10376 19320 10382 19372
rect 10520 19369 10548 19400
rect 10594 19388 10600 19440
rect 10652 19428 10658 19440
rect 10778 19428 10784 19440
rect 10652 19400 10784 19428
rect 10652 19388 10658 19400
rect 10778 19388 10784 19400
rect 10836 19388 10842 19440
rect 10962 19388 10968 19440
rect 11020 19428 11026 19440
rect 11609 19431 11667 19437
rect 11609 19428 11621 19431
rect 11020 19400 11621 19428
rect 11020 19388 11026 19400
rect 11609 19397 11621 19400
rect 11655 19397 11667 19431
rect 11609 19391 11667 19397
rect 11793 19431 11851 19437
rect 11793 19397 11805 19431
rect 11839 19428 11851 19431
rect 11974 19428 11980 19440
rect 11839 19400 11980 19428
rect 11839 19397 11851 19400
rect 11793 19391 11851 19397
rect 11974 19388 11980 19400
rect 12032 19388 12038 19440
rect 12342 19388 12348 19440
rect 12400 19428 12406 19440
rect 12621 19431 12679 19437
rect 12621 19428 12633 19431
rect 12400 19400 12633 19428
rect 12400 19388 12406 19400
rect 12621 19397 12633 19400
rect 12667 19397 12679 19431
rect 14185 19431 14243 19437
rect 14185 19428 14197 19431
rect 12621 19391 12679 19397
rect 13280 19400 14197 19428
rect 10505 19363 10563 19369
rect 10505 19329 10517 19363
rect 10551 19329 10563 19363
rect 13280 19360 13308 19400
rect 14185 19397 14197 19400
rect 14231 19397 14243 19431
rect 14185 19391 14243 19397
rect 19153 19431 19211 19437
rect 19153 19397 19165 19431
rect 19199 19428 19211 19431
rect 19794 19428 19800 19440
rect 19199 19400 19800 19428
rect 19199 19397 19211 19400
rect 19153 19391 19211 19397
rect 19794 19388 19800 19400
rect 19852 19388 19858 19440
rect 13446 19360 13452 19372
rect 10505 19323 10563 19329
rect 12268 19332 13308 19360
rect 13407 19332 13452 19360
rect 12268 19304 12296 19332
rect 13446 19320 13452 19332
rect 13504 19320 13510 19372
rect 13630 19360 13636 19372
rect 13591 19332 13636 19360
rect 13630 19320 13636 19332
rect 13688 19320 13694 19372
rect 13725 19363 13783 19369
rect 13725 19329 13737 19363
rect 13771 19329 13783 19363
rect 13725 19323 13783 19329
rect 10594 19292 10600 19304
rect 10555 19264 10600 19292
rect 10594 19252 10600 19264
rect 10652 19252 10658 19304
rect 12250 19292 12256 19304
rect 12211 19264 12256 19292
rect 12250 19252 12256 19264
rect 12308 19252 12314 19304
rect 12710 19292 12716 19304
rect 12406 19264 12716 19292
rect 12406 19236 12434 19264
rect 12710 19252 12716 19264
rect 12768 19252 12774 19304
rect 13170 19292 13176 19304
rect 12820 19264 13176 19292
rect 10778 19184 10784 19236
rect 10836 19224 10842 19236
rect 12406 19224 12440 19236
rect 10836 19196 12440 19224
rect 10836 19184 10842 19196
rect 12434 19184 12440 19196
rect 12492 19184 12498 19236
rect 12820 19233 12848 19264
rect 13170 19252 13176 19264
rect 13228 19292 13234 19304
rect 13740 19292 13768 19323
rect 13814 19320 13820 19372
rect 13872 19360 13878 19372
rect 14369 19363 14427 19369
rect 14369 19360 14381 19363
rect 13872 19332 14381 19360
rect 13872 19320 13878 19332
rect 14369 19329 14381 19332
rect 14415 19329 14427 19363
rect 14369 19323 14427 19329
rect 14461 19363 14519 19369
rect 14461 19329 14473 19363
rect 14507 19329 14519 19363
rect 15378 19360 15384 19372
rect 15339 19332 15384 19360
rect 14461 19323 14519 19329
rect 13228 19264 13768 19292
rect 13228 19252 13234 19264
rect 12805 19227 12863 19233
rect 12805 19193 12817 19227
rect 12851 19193 12863 19227
rect 14476 19224 14504 19323
rect 15378 19320 15384 19332
rect 15436 19320 15442 19372
rect 16942 19360 16948 19372
rect 16903 19332 16948 19360
rect 16942 19320 16948 19332
rect 17000 19320 17006 19372
rect 17218 19369 17224 19372
rect 17212 19323 17224 19369
rect 17276 19360 17282 19372
rect 17276 19332 17312 19360
rect 17218 19320 17224 19323
rect 17276 19320 17282 19332
rect 18782 19320 18788 19372
rect 18840 19360 18846 19372
rect 18877 19363 18935 19369
rect 18877 19360 18889 19363
rect 18840 19332 18889 19360
rect 18840 19320 18846 19332
rect 18877 19329 18889 19332
rect 18923 19329 18935 19363
rect 18877 19323 18935 19329
rect 19061 19363 19119 19369
rect 19061 19329 19073 19363
rect 19107 19329 19119 19363
rect 19061 19323 19119 19329
rect 15654 19292 15660 19304
rect 15615 19264 15660 19292
rect 15654 19252 15660 19264
rect 15712 19252 15718 19304
rect 19076 19292 19104 19323
rect 19242 19320 19248 19372
rect 19300 19360 19306 19372
rect 20088 19369 20116 19468
rect 20346 19456 20352 19468
rect 20404 19456 20410 19508
rect 20441 19499 20499 19505
rect 20441 19465 20453 19499
rect 20487 19496 20499 19499
rect 21082 19496 21088 19508
rect 20487 19468 21088 19496
rect 20487 19465 20499 19468
rect 20441 19459 20499 19465
rect 21082 19456 21088 19468
rect 21140 19456 21146 19508
rect 22738 19456 22744 19508
rect 22796 19496 22802 19508
rect 23017 19499 23075 19505
rect 23017 19496 23029 19499
rect 22796 19468 23029 19496
rect 22796 19456 22802 19468
rect 23017 19465 23029 19468
rect 23063 19465 23075 19499
rect 25590 19496 25596 19508
rect 25551 19468 25596 19496
rect 23017 19459 23075 19465
rect 25590 19456 25596 19468
rect 25648 19456 25654 19508
rect 25700 19468 25912 19496
rect 20165 19431 20223 19437
rect 20165 19397 20177 19431
rect 20211 19428 20223 19431
rect 20898 19428 20904 19440
rect 20211 19400 20904 19428
rect 20211 19397 20223 19400
rect 20165 19391 20223 19397
rect 20898 19388 20904 19400
rect 20956 19388 20962 19440
rect 22646 19428 22652 19440
rect 21376 19400 22652 19428
rect 19889 19363 19947 19369
rect 19300 19332 19840 19360
rect 19300 19320 19306 19332
rect 19812 19304 19840 19332
rect 19889 19329 19901 19363
rect 19935 19360 19947 19363
rect 20073 19363 20131 19369
rect 19935 19332 20024 19360
rect 19935 19329 19947 19332
rect 19889 19323 19947 19329
rect 19150 19292 19156 19304
rect 19076 19264 19156 19292
rect 19150 19252 19156 19264
rect 19208 19252 19214 19304
rect 19794 19252 19800 19304
rect 19852 19252 19858 19304
rect 19996 19284 20024 19332
rect 20073 19329 20085 19363
rect 20119 19329 20131 19363
rect 20073 19323 20131 19329
rect 20257 19363 20315 19369
rect 20257 19329 20269 19363
rect 20303 19329 20315 19363
rect 20257 19323 20315 19329
rect 19904 19256 20024 19284
rect 16758 19224 16764 19236
rect 12805 19187 12863 19193
rect 12912 19196 14504 19224
rect 14568 19196 16764 19224
rect 12618 19156 12624 19168
rect 12531 19128 12624 19156
rect 12618 19116 12624 19128
rect 12676 19156 12682 19168
rect 12912 19156 12940 19196
rect 12676 19128 12940 19156
rect 12676 19116 12682 19128
rect 12986 19116 12992 19168
rect 13044 19156 13050 19168
rect 13265 19159 13323 19165
rect 13265 19156 13277 19159
rect 13044 19128 13277 19156
rect 13044 19116 13050 19128
rect 13265 19125 13277 19128
rect 13311 19125 13323 19159
rect 13265 19119 13323 19125
rect 13354 19116 13360 19168
rect 13412 19156 13418 19168
rect 14568 19156 14596 19196
rect 16758 19184 16764 19196
rect 16816 19184 16822 19236
rect 15010 19156 15016 19168
rect 13412 19128 14596 19156
rect 14971 19128 15016 19156
rect 13412 19116 13418 19128
rect 15010 19116 15016 19128
rect 15068 19116 15074 19168
rect 15102 19116 15108 19168
rect 15160 19156 15166 19168
rect 19904 19156 19932 19256
rect 20272 19224 20300 19323
rect 20530 19320 20536 19372
rect 20588 19360 20594 19372
rect 20993 19363 21051 19369
rect 20993 19360 21005 19363
rect 20588 19332 21005 19360
rect 20588 19320 20594 19332
rect 20993 19329 21005 19332
rect 21039 19329 21051 19363
rect 21376 19360 21404 19400
rect 22646 19388 22652 19400
rect 22704 19388 22710 19440
rect 20993 19323 21051 19329
rect 21284 19332 21404 19360
rect 22281 19363 22339 19369
rect 20346 19252 20352 19304
rect 20404 19292 20410 19304
rect 21284 19292 21312 19332
rect 22281 19329 22293 19363
rect 22327 19360 22339 19363
rect 23750 19360 23756 19372
rect 22327 19332 23756 19360
rect 22327 19329 22339 19332
rect 22281 19323 22339 19329
rect 23750 19320 23756 19332
rect 23808 19320 23814 19372
rect 23842 19320 23848 19372
rect 23900 19360 23906 19372
rect 24029 19363 24087 19369
rect 24029 19360 24041 19363
rect 23900 19332 24041 19360
rect 23900 19320 23906 19332
rect 24029 19329 24041 19332
rect 24075 19360 24087 19363
rect 25498 19360 25504 19372
rect 24075 19332 25504 19360
rect 24075 19329 24087 19332
rect 24029 19323 24087 19329
rect 25498 19320 25504 19332
rect 25556 19320 25562 19372
rect 25590 19320 25596 19372
rect 25648 19360 25654 19372
rect 25700 19360 25728 19468
rect 25884 19437 25912 19468
rect 26234 19456 26240 19508
rect 26292 19496 26298 19508
rect 29914 19496 29920 19508
rect 26292 19468 29920 19496
rect 26292 19456 26298 19468
rect 25869 19431 25927 19437
rect 25869 19397 25881 19431
rect 25915 19397 25927 19431
rect 25869 19391 25927 19397
rect 26099 19431 26157 19437
rect 26099 19397 26111 19431
rect 26145 19428 26157 19431
rect 27338 19428 27344 19440
rect 26145 19400 27344 19428
rect 26145 19397 26157 19400
rect 26099 19391 26157 19397
rect 27338 19388 27344 19400
rect 27396 19388 27402 19440
rect 29638 19428 29644 19440
rect 29599 19400 29644 19428
rect 29638 19388 29644 19400
rect 29696 19388 29702 19440
rect 29748 19437 29776 19468
rect 29914 19456 29920 19468
rect 29972 19456 29978 19508
rect 33870 19496 33876 19508
rect 33831 19468 33876 19496
rect 33870 19456 33876 19468
rect 33928 19456 33934 19508
rect 34974 19456 34980 19508
rect 35032 19496 35038 19508
rect 35253 19499 35311 19505
rect 35253 19496 35265 19499
rect 35032 19468 35265 19496
rect 35032 19456 35038 19468
rect 35253 19465 35265 19468
rect 35299 19465 35311 19499
rect 35253 19459 35311 19465
rect 29733 19431 29791 19437
rect 29733 19397 29745 19431
rect 29779 19397 29791 19431
rect 29733 19391 29791 19397
rect 30558 19388 30564 19440
rect 30616 19428 30622 19440
rect 30653 19431 30711 19437
rect 30653 19428 30665 19431
rect 30616 19400 30665 19428
rect 30616 19388 30622 19400
rect 30653 19397 30665 19400
rect 30699 19397 30711 19431
rect 30653 19391 30711 19397
rect 30837 19431 30895 19437
rect 30837 19397 30849 19431
rect 30883 19428 30895 19431
rect 31110 19428 31116 19440
rect 30883 19400 31116 19428
rect 30883 19397 30895 19400
rect 30837 19391 30895 19397
rect 31110 19388 31116 19400
rect 31168 19388 31174 19440
rect 32582 19388 32588 19440
rect 32640 19428 32646 19440
rect 32858 19428 32864 19440
rect 32640 19400 32864 19428
rect 32640 19388 32646 19400
rect 32858 19388 32864 19400
rect 32916 19428 32922 19440
rect 35342 19428 35348 19440
rect 32916 19400 35348 19428
rect 32916 19388 32922 19400
rect 25648 19332 25728 19360
rect 25648 19320 25654 19332
rect 25774 19320 25780 19372
rect 25832 19360 25838 19372
rect 25961 19363 26019 19369
rect 25832 19332 25877 19360
rect 25832 19320 25838 19332
rect 25961 19329 25973 19363
rect 26007 19360 26019 19363
rect 26234 19360 26240 19372
rect 26007 19332 26041 19360
rect 26195 19332 26240 19360
rect 26007 19329 26019 19332
rect 25961 19323 26019 19329
rect 20404 19264 21312 19292
rect 20404 19252 20410 19264
rect 21910 19252 21916 19304
rect 21968 19292 21974 19304
rect 22005 19295 22063 19301
rect 22005 19292 22017 19295
rect 21968 19264 22017 19292
rect 21968 19252 21974 19264
rect 22005 19261 22017 19264
rect 22051 19261 22063 19295
rect 22005 19255 22063 19261
rect 24305 19295 24363 19301
rect 24305 19261 24317 19295
rect 24351 19292 24363 19295
rect 24486 19292 24492 19304
rect 24351 19264 24492 19292
rect 24351 19261 24363 19264
rect 24305 19255 24363 19261
rect 24486 19252 24492 19264
rect 24544 19292 24550 19304
rect 25976 19292 26004 19323
rect 26234 19320 26240 19332
rect 26292 19320 26298 19372
rect 27525 19363 27583 19369
rect 27525 19329 27537 19363
rect 27571 19360 27583 19363
rect 28442 19360 28448 19372
rect 27571 19332 28448 19360
rect 27571 19329 27583 19332
rect 27525 19323 27583 19329
rect 28442 19320 28448 19332
rect 28500 19320 28506 19372
rect 28537 19363 28595 19369
rect 28537 19329 28549 19363
rect 28583 19360 28595 19363
rect 28994 19360 29000 19372
rect 28583 19332 29000 19360
rect 28583 19329 28595 19332
rect 28537 19323 28595 19329
rect 28994 19320 29000 19332
rect 29052 19320 29058 19372
rect 29546 19360 29552 19372
rect 29507 19332 29552 19360
rect 29546 19320 29552 19332
rect 29604 19320 29610 19372
rect 29851 19363 29909 19369
rect 29851 19360 29863 19363
rect 29748 19332 29863 19360
rect 26050 19292 26056 19304
rect 24544 19264 25912 19292
rect 25976 19264 26056 19292
rect 24544 19252 24550 19264
rect 20530 19224 20536 19236
rect 20272 19196 20536 19224
rect 20530 19184 20536 19196
rect 20588 19184 20594 19236
rect 20990 19184 20996 19236
rect 21048 19224 21054 19236
rect 21928 19224 21956 19252
rect 21048 19196 21956 19224
rect 21048 19184 21054 19196
rect 23566 19184 23572 19236
rect 23624 19224 23630 19236
rect 25774 19224 25780 19236
rect 23624 19196 25780 19224
rect 23624 19184 23630 19196
rect 25774 19184 25780 19196
rect 25832 19184 25838 19236
rect 25884 19224 25912 19264
rect 26050 19252 26056 19264
rect 26108 19252 26114 19304
rect 27801 19295 27859 19301
rect 27801 19292 27813 19295
rect 26160 19264 27813 19292
rect 26160 19224 26188 19264
rect 27801 19261 27813 19264
rect 27847 19261 27859 19295
rect 27801 19255 27859 19261
rect 28629 19295 28687 19301
rect 28629 19261 28641 19295
rect 28675 19261 28687 19295
rect 28629 19255 28687 19261
rect 28905 19295 28963 19301
rect 28905 19261 28917 19295
rect 28951 19292 28963 19295
rect 29748 19292 29776 19332
rect 29851 19329 29863 19332
rect 29897 19329 29909 19363
rect 32122 19360 32128 19372
rect 32083 19332 32128 19360
rect 29851 19323 29909 19329
rect 32122 19320 32128 19332
rect 32180 19320 32186 19372
rect 32309 19363 32367 19369
rect 32309 19329 32321 19363
rect 32355 19329 32367 19363
rect 32309 19323 32367 19329
rect 28951 19264 29776 19292
rect 30009 19295 30067 19301
rect 28951 19261 28963 19264
rect 28905 19255 28963 19261
rect 30009 19261 30021 19295
rect 30055 19292 30067 19295
rect 30190 19292 30196 19304
rect 30055 19264 30196 19292
rect 30055 19261 30067 19264
rect 30009 19255 30067 19261
rect 25884 19196 26188 19224
rect 27617 19227 27675 19233
rect 27617 19193 27629 19227
rect 27663 19224 27675 19227
rect 27890 19224 27896 19236
rect 27663 19196 27896 19224
rect 27663 19193 27675 19196
rect 27617 19187 27675 19193
rect 27890 19184 27896 19196
rect 27948 19184 27954 19236
rect 20254 19156 20260 19168
rect 15160 19128 20260 19156
rect 15160 19116 15166 19128
rect 20254 19116 20260 19128
rect 20312 19116 20318 19168
rect 20806 19116 20812 19168
rect 20864 19156 20870 19168
rect 21085 19159 21143 19165
rect 21085 19156 21097 19159
rect 20864 19128 21097 19156
rect 20864 19116 20870 19128
rect 21085 19125 21097 19128
rect 21131 19156 21143 19159
rect 23290 19156 23296 19168
rect 21131 19128 23296 19156
rect 21131 19125 21143 19128
rect 21085 19119 21143 19125
rect 23290 19116 23296 19128
rect 23348 19116 23354 19168
rect 25682 19116 25688 19168
rect 25740 19156 25746 19168
rect 26050 19156 26056 19168
rect 25740 19128 26056 19156
rect 25740 19116 25746 19128
rect 26050 19116 26056 19128
rect 26108 19116 26114 19168
rect 26234 19116 26240 19168
rect 26292 19156 26298 19168
rect 27709 19159 27767 19165
rect 27709 19156 27721 19159
rect 26292 19128 27721 19156
rect 26292 19116 26298 19128
rect 27709 19125 27721 19128
rect 27755 19125 27767 19159
rect 28644 19156 28672 19255
rect 30190 19252 30196 19264
rect 30248 19252 30254 19304
rect 31754 19252 31760 19304
rect 31812 19292 31818 19304
rect 32324 19292 32352 19323
rect 32674 19320 32680 19372
rect 32732 19360 32738 19372
rect 33244 19369 33272 19400
rect 35342 19388 35348 19400
rect 35400 19388 35406 19440
rect 33009 19363 33067 19369
rect 33009 19360 33021 19363
rect 32732 19332 33021 19360
rect 32732 19320 32738 19332
rect 33009 19329 33021 19332
rect 33055 19329 33067 19363
rect 33009 19323 33067 19329
rect 33137 19363 33195 19369
rect 33137 19329 33149 19363
rect 33183 19329 33195 19363
rect 33137 19323 33195 19329
rect 33229 19363 33287 19369
rect 33229 19329 33241 19363
rect 33275 19329 33287 19363
rect 34054 19360 34060 19372
rect 34015 19332 34060 19360
rect 33229 19323 33287 19329
rect 31812 19264 32352 19292
rect 33152 19292 33180 19323
rect 34054 19320 34060 19332
rect 34112 19320 34118 19372
rect 34146 19320 34152 19372
rect 34204 19360 34210 19372
rect 34425 19363 34483 19369
rect 34204 19332 34249 19360
rect 34204 19320 34210 19332
rect 34425 19329 34437 19363
rect 34471 19329 34483 19363
rect 34425 19323 34483 19329
rect 34440 19292 34468 19323
rect 34606 19320 34612 19372
rect 34664 19360 34670 19372
rect 34885 19363 34943 19369
rect 34885 19360 34897 19363
rect 34664 19332 34897 19360
rect 34664 19320 34670 19332
rect 34885 19329 34897 19332
rect 34931 19329 34943 19363
rect 34885 19323 34943 19329
rect 33152 19264 33272 19292
rect 31812 19252 31818 19264
rect 28718 19184 28724 19236
rect 28776 19224 28782 19236
rect 32398 19224 32404 19236
rect 28776 19196 32404 19224
rect 28776 19184 28782 19196
rect 32398 19184 32404 19196
rect 32456 19184 32462 19236
rect 33134 19184 33140 19236
rect 33192 19224 33198 19236
rect 33244 19224 33272 19264
rect 33192 19196 33272 19224
rect 33980 19264 34468 19292
rect 33192 19184 33198 19196
rect 33980 19168 34008 19264
rect 34698 19252 34704 19304
rect 34756 19292 34762 19304
rect 34977 19295 35035 19301
rect 34977 19292 34989 19295
rect 34756 19264 34989 19292
rect 34756 19252 34762 19264
rect 34977 19261 34989 19264
rect 35023 19261 35035 19295
rect 34977 19255 35035 19261
rect 34333 19227 34391 19233
rect 34333 19193 34345 19227
rect 34379 19224 34391 19227
rect 34790 19224 34796 19236
rect 34379 19196 34796 19224
rect 34379 19193 34391 19196
rect 34333 19187 34391 19193
rect 34790 19184 34796 19196
rect 34848 19184 34854 19236
rect 29086 19156 29092 19168
rect 28644 19128 29092 19156
rect 27709 19119 27767 19125
rect 29086 19116 29092 19128
rect 29144 19116 29150 19168
rect 29362 19156 29368 19168
rect 29323 19128 29368 19156
rect 29362 19116 29368 19128
rect 29420 19116 29426 19168
rect 31021 19159 31079 19165
rect 31021 19125 31033 19159
rect 31067 19156 31079 19159
rect 31110 19156 31116 19168
rect 31067 19128 31116 19156
rect 31067 19125 31079 19128
rect 31021 19119 31079 19125
rect 31110 19116 31116 19128
rect 31168 19116 31174 19168
rect 31294 19116 31300 19168
rect 31352 19156 31358 19168
rect 32125 19159 32183 19165
rect 32125 19156 32137 19159
rect 31352 19128 32137 19156
rect 31352 19116 31358 19128
rect 32125 19125 32137 19128
rect 32171 19125 32183 19159
rect 32125 19119 32183 19125
rect 33413 19159 33471 19165
rect 33413 19125 33425 19159
rect 33459 19156 33471 19159
rect 33962 19156 33968 19168
rect 33459 19128 33968 19156
rect 33459 19125 33471 19128
rect 33413 19119 33471 19125
rect 33962 19116 33968 19128
rect 34020 19116 34026 19168
rect 35069 19159 35127 19165
rect 35069 19125 35081 19159
rect 35115 19156 35127 19159
rect 35526 19156 35532 19168
rect 35115 19128 35532 19156
rect 35115 19125 35127 19128
rect 35069 19119 35127 19125
rect 35526 19116 35532 19128
rect 35584 19116 35590 19168
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 8018 18912 8024 18964
rect 8076 18952 8082 18964
rect 8113 18955 8171 18961
rect 8113 18952 8125 18955
rect 8076 18924 8125 18952
rect 8076 18912 8082 18924
rect 8113 18921 8125 18924
rect 8159 18921 8171 18955
rect 8113 18915 8171 18921
rect 9585 18955 9643 18961
rect 9585 18921 9597 18955
rect 9631 18952 9643 18955
rect 10318 18952 10324 18964
rect 9631 18924 10324 18952
rect 9631 18921 9643 18924
rect 9585 18915 9643 18921
rect 10318 18912 10324 18924
rect 10376 18912 10382 18964
rect 10594 18912 10600 18964
rect 10652 18952 10658 18964
rect 11241 18955 11299 18961
rect 11241 18952 11253 18955
rect 10652 18924 11253 18952
rect 10652 18912 10658 18924
rect 11241 18921 11253 18924
rect 11287 18921 11299 18955
rect 11241 18915 11299 18921
rect 13541 18955 13599 18961
rect 13541 18921 13553 18955
rect 13587 18952 13599 18955
rect 13814 18952 13820 18964
rect 13587 18924 13820 18952
rect 13587 18921 13599 18924
rect 13541 18915 13599 18921
rect 13814 18912 13820 18924
rect 13872 18912 13878 18964
rect 13906 18912 13912 18964
rect 13964 18952 13970 18964
rect 15102 18952 15108 18964
rect 13964 18924 15108 18952
rect 13964 18912 13970 18924
rect 15102 18912 15108 18924
rect 15160 18912 15166 18964
rect 15378 18912 15384 18964
rect 15436 18952 15442 18964
rect 15749 18955 15807 18961
rect 15749 18952 15761 18955
rect 15436 18924 15761 18952
rect 15436 18912 15442 18924
rect 15749 18921 15761 18924
rect 15795 18921 15807 18955
rect 15749 18915 15807 18921
rect 15764 18884 15792 18915
rect 16758 18912 16764 18964
rect 16816 18952 16822 18964
rect 16816 18924 17172 18952
rect 16816 18912 16822 18924
rect 15764 18856 17080 18884
rect 10226 18816 10232 18828
rect 10187 18788 10232 18816
rect 10226 18776 10232 18788
rect 10284 18776 10290 18828
rect 11609 18819 11667 18825
rect 11609 18816 11621 18819
rect 10336 18788 11621 18816
rect 8294 18748 8300 18760
rect 8255 18720 8300 18748
rect 8294 18708 8300 18720
rect 8352 18708 8358 18760
rect 9493 18751 9551 18757
rect 9493 18717 9505 18751
rect 9539 18717 9551 18751
rect 9674 18748 9680 18760
rect 9635 18720 9680 18748
rect 9493 18711 9551 18717
rect 9508 18680 9536 18711
rect 9674 18708 9680 18720
rect 9732 18708 9738 18760
rect 10336 18757 10364 18788
rect 11609 18785 11621 18788
rect 11655 18785 11667 18819
rect 16942 18816 16948 18828
rect 11609 18779 11667 18785
rect 15672 18788 16948 18816
rect 10321 18751 10379 18757
rect 10321 18717 10333 18751
rect 10367 18717 10379 18751
rect 10321 18711 10379 18717
rect 10410 18708 10416 18760
rect 10468 18748 10474 18760
rect 11149 18751 11207 18757
rect 11149 18748 11161 18751
rect 10468 18720 11161 18748
rect 10468 18708 10474 18720
rect 11149 18717 11161 18720
rect 11195 18717 11207 18751
rect 11149 18711 11207 18717
rect 11882 18708 11888 18760
rect 11940 18748 11946 18760
rect 12161 18751 12219 18757
rect 12161 18748 12173 18751
rect 11940 18720 12173 18748
rect 11940 18708 11946 18720
rect 12161 18717 12173 18720
rect 12207 18717 12219 18751
rect 14366 18748 14372 18760
rect 14279 18720 14372 18748
rect 12161 18711 12219 18717
rect 14366 18708 14372 18720
rect 14424 18748 14430 18760
rect 15672 18748 15700 18788
rect 16942 18776 16948 18788
rect 17000 18776 17006 18828
rect 16390 18748 16396 18760
rect 14424 18720 15700 18748
rect 16351 18720 16396 18748
rect 14424 18708 14430 18720
rect 16390 18708 16396 18720
rect 16448 18708 16454 18760
rect 16853 18751 16911 18757
rect 16853 18717 16865 18751
rect 16899 18748 16911 18751
rect 17052 18748 17080 18856
rect 16899 18720 17080 18748
rect 17144 18748 17172 18924
rect 19334 18912 19340 18964
rect 19392 18952 19398 18964
rect 20993 18955 21051 18961
rect 20993 18952 21005 18955
rect 19392 18924 21005 18952
rect 19392 18912 19398 18924
rect 20993 18921 21005 18924
rect 21039 18921 21051 18955
rect 20993 18915 21051 18921
rect 22002 18912 22008 18964
rect 22060 18912 22066 18964
rect 23566 18912 23572 18964
rect 23624 18952 23630 18964
rect 23661 18955 23719 18961
rect 23661 18952 23673 18955
rect 23624 18924 23673 18952
rect 23624 18912 23630 18924
rect 23661 18921 23673 18924
rect 23707 18921 23719 18955
rect 23842 18952 23848 18964
rect 23803 18924 23848 18952
rect 23661 18915 23719 18921
rect 23842 18912 23848 18924
rect 23900 18912 23906 18964
rect 24854 18912 24860 18964
rect 24912 18952 24918 18964
rect 26145 18955 26203 18961
rect 26145 18952 26157 18955
rect 24912 18924 26157 18952
rect 24912 18912 24918 18924
rect 26145 18921 26157 18924
rect 26191 18921 26203 18955
rect 26145 18915 26203 18921
rect 27890 18912 27896 18964
rect 27948 18952 27954 18964
rect 28169 18955 28227 18961
rect 28169 18952 28181 18955
rect 27948 18924 28181 18952
rect 27948 18912 27954 18924
rect 28169 18921 28181 18924
rect 28215 18921 28227 18955
rect 28169 18915 28227 18921
rect 29270 18912 29276 18964
rect 29328 18952 29334 18964
rect 29549 18955 29607 18961
rect 29549 18952 29561 18955
rect 29328 18924 29561 18952
rect 29328 18912 29334 18924
rect 29549 18921 29561 18924
rect 29595 18921 29607 18955
rect 29549 18915 29607 18921
rect 29656 18924 30144 18952
rect 17954 18844 17960 18896
rect 18012 18884 18018 18896
rect 18012 18856 18092 18884
rect 18012 18844 18018 18856
rect 18064 18757 18092 18856
rect 18690 18844 18696 18896
rect 18748 18884 18754 18896
rect 22020 18884 22048 18912
rect 18748 18856 22048 18884
rect 18748 18844 18754 18856
rect 23290 18844 23296 18896
rect 23348 18884 23354 18896
rect 24670 18884 24676 18896
rect 23348 18856 24676 18884
rect 23348 18844 23354 18856
rect 18414 18776 18420 18828
rect 18472 18816 18478 18828
rect 20898 18816 20904 18828
rect 18472 18788 20904 18816
rect 18472 18776 18478 18788
rect 20898 18776 20904 18788
rect 20956 18776 20962 18828
rect 23771 18825 23799 18856
rect 24670 18844 24676 18856
rect 24728 18844 24734 18896
rect 24765 18887 24823 18893
rect 24765 18853 24777 18887
rect 24811 18884 24823 18887
rect 29362 18884 29368 18896
rect 24811 18856 29368 18884
rect 24811 18853 24823 18856
rect 24765 18847 24823 18853
rect 29362 18844 29368 18856
rect 29420 18844 29426 18896
rect 23753 18819 23811 18825
rect 23753 18785 23765 18819
rect 23799 18785 23811 18819
rect 23753 18779 23811 18785
rect 24302 18776 24308 18828
rect 24360 18816 24366 18828
rect 29656 18816 29684 18924
rect 24360 18788 29684 18816
rect 30116 18816 30144 18924
rect 30466 18912 30472 18964
rect 30524 18952 30530 18964
rect 30653 18955 30711 18961
rect 30653 18952 30665 18955
rect 30524 18924 30665 18952
rect 30524 18912 30530 18924
rect 30653 18921 30665 18924
rect 30699 18921 30711 18955
rect 30653 18915 30711 18921
rect 31754 18912 31760 18964
rect 31812 18952 31818 18964
rect 31812 18924 31857 18952
rect 31812 18912 31818 18924
rect 34054 18844 34060 18896
rect 34112 18884 34118 18896
rect 35253 18887 35311 18893
rect 35253 18884 35265 18887
rect 34112 18856 35265 18884
rect 34112 18844 34118 18856
rect 35253 18853 35265 18856
rect 35299 18853 35311 18887
rect 35253 18847 35311 18853
rect 34514 18816 34520 18828
rect 30116 18788 34520 18816
rect 24360 18776 24366 18788
rect 34514 18776 34520 18788
rect 34572 18776 34578 18828
rect 34974 18816 34980 18828
rect 34935 18788 34980 18816
rect 34974 18776 34980 18788
rect 35032 18776 35038 18828
rect 17865 18751 17923 18757
rect 17865 18748 17877 18751
rect 17144 18720 17877 18748
rect 16899 18717 16911 18720
rect 16853 18711 16911 18717
rect 17865 18717 17877 18720
rect 17911 18717 17923 18751
rect 17865 18711 17923 18717
rect 18049 18751 18107 18757
rect 18049 18717 18061 18751
rect 18095 18717 18107 18751
rect 18230 18748 18236 18760
rect 18191 18720 18236 18748
rect 18049 18711 18107 18717
rect 18230 18708 18236 18720
rect 18288 18708 18294 18760
rect 19702 18748 19708 18760
rect 19663 18720 19708 18748
rect 19702 18708 19708 18720
rect 19760 18708 19766 18760
rect 21910 18748 21916 18760
rect 21871 18720 21916 18748
rect 21910 18708 21916 18720
rect 21968 18708 21974 18760
rect 22189 18751 22247 18757
rect 22189 18717 22201 18751
rect 22235 18748 22247 18751
rect 23106 18748 23112 18760
rect 22235 18720 23112 18748
rect 22235 18717 22247 18720
rect 22189 18711 22247 18717
rect 23106 18708 23112 18720
rect 23164 18708 23170 18760
rect 23569 18751 23627 18757
rect 23569 18717 23581 18751
rect 23615 18748 23627 18751
rect 24486 18748 24492 18760
rect 23615 18720 24492 18748
rect 23615 18717 23627 18720
rect 23569 18711 23627 18717
rect 24486 18708 24492 18720
rect 24544 18748 24550 18760
rect 24581 18751 24639 18757
rect 24581 18748 24593 18751
rect 24544 18720 24593 18748
rect 24544 18708 24550 18720
rect 24581 18717 24593 18720
rect 24627 18717 24639 18751
rect 24581 18711 24639 18717
rect 24673 18751 24731 18757
rect 24673 18717 24685 18751
rect 24719 18717 24731 18751
rect 24673 18711 24731 18717
rect 24857 18751 24915 18757
rect 24857 18717 24869 18751
rect 24903 18717 24915 18751
rect 25038 18748 25044 18760
rect 24999 18720 25044 18748
rect 24857 18711 24915 18717
rect 9766 18680 9772 18692
rect 9508 18652 9772 18680
rect 9766 18640 9772 18652
rect 9824 18640 9830 18692
rect 12428 18683 12486 18689
rect 12428 18649 12440 18683
rect 12474 18680 12486 18683
rect 12710 18680 12716 18692
rect 12474 18652 12716 18680
rect 12474 18649 12486 18652
rect 12428 18643 12486 18649
rect 12710 18640 12716 18652
rect 12768 18640 12774 18692
rect 14636 18683 14694 18689
rect 14636 18649 14648 18683
rect 14682 18680 14694 18683
rect 16209 18683 16267 18689
rect 16209 18680 16221 18683
rect 14682 18652 16221 18680
rect 14682 18649 14694 18652
rect 14636 18643 14694 18649
rect 16209 18649 16221 18652
rect 16255 18649 16267 18683
rect 16209 18643 16267 18649
rect 16298 18640 16304 18692
rect 16356 18680 16362 18692
rect 16485 18683 16543 18689
rect 16485 18680 16497 18683
rect 16356 18652 16497 18680
rect 16356 18640 16362 18652
rect 16485 18649 16497 18652
rect 16531 18649 16543 18683
rect 16485 18643 16543 18649
rect 16574 18640 16580 18692
rect 16632 18680 16638 18692
rect 16758 18689 16764 18692
rect 16715 18683 16764 18689
rect 16632 18652 16677 18680
rect 16632 18640 16638 18652
rect 16715 18649 16727 18683
rect 16761 18649 16764 18683
rect 16715 18643 16764 18649
rect 16758 18640 16764 18643
rect 16816 18640 16822 18692
rect 18138 18640 18144 18692
rect 18196 18680 18202 18692
rect 23385 18683 23443 18689
rect 18196 18652 18241 18680
rect 18196 18640 18202 18652
rect 23385 18649 23397 18683
rect 23431 18680 23443 18683
rect 24118 18680 24124 18692
rect 23431 18652 24124 18680
rect 23431 18649 23443 18652
rect 23385 18643 23443 18649
rect 24118 18640 24124 18652
rect 24176 18640 24182 18692
rect 10689 18615 10747 18621
rect 10689 18581 10701 18615
rect 10735 18612 10747 18615
rect 11238 18612 11244 18624
rect 10735 18584 11244 18612
rect 10735 18581 10747 18584
rect 10689 18575 10747 18581
rect 11238 18572 11244 18584
rect 11296 18572 11302 18624
rect 17954 18572 17960 18624
rect 18012 18612 18018 18624
rect 18417 18615 18475 18621
rect 18417 18612 18429 18615
rect 18012 18584 18429 18612
rect 18012 18572 18018 18584
rect 18417 18581 18429 18584
rect 18463 18581 18475 18615
rect 18417 18575 18475 18581
rect 18966 18572 18972 18624
rect 19024 18612 19030 18624
rect 21818 18612 21824 18624
rect 19024 18584 21824 18612
rect 19024 18572 19030 18584
rect 21818 18572 21824 18584
rect 21876 18572 21882 18624
rect 21910 18572 21916 18624
rect 21968 18612 21974 18624
rect 22738 18612 22744 18624
rect 21968 18584 22744 18612
rect 21968 18572 21974 18584
rect 22738 18572 22744 18584
rect 22796 18572 22802 18624
rect 22925 18615 22983 18621
rect 22925 18581 22937 18615
rect 22971 18612 22983 18615
rect 23290 18612 23296 18624
rect 22971 18584 23296 18612
rect 22971 18581 22983 18584
rect 22925 18575 22983 18581
rect 23290 18572 23296 18584
rect 23348 18572 23354 18624
rect 23566 18572 23572 18624
rect 23624 18612 23630 18624
rect 24397 18615 24455 18621
rect 24397 18612 24409 18615
rect 23624 18584 24409 18612
rect 23624 18572 23630 18584
rect 24397 18581 24409 18584
rect 24443 18581 24455 18615
rect 24688 18612 24716 18711
rect 24872 18680 24900 18711
rect 25038 18708 25044 18720
rect 25096 18708 25102 18760
rect 25498 18748 25504 18760
rect 25459 18720 25504 18748
rect 25498 18708 25504 18720
rect 25556 18708 25562 18760
rect 25866 18748 25872 18760
rect 25827 18720 25872 18748
rect 25866 18708 25872 18720
rect 25924 18708 25930 18760
rect 25961 18751 26019 18757
rect 25961 18717 25973 18751
rect 26007 18748 26019 18751
rect 26326 18748 26332 18760
rect 26007 18720 26332 18748
rect 26007 18717 26019 18720
rect 25961 18711 26019 18717
rect 26326 18708 26332 18720
rect 26384 18748 26390 18760
rect 26605 18751 26663 18757
rect 26605 18748 26617 18751
rect 26384 18720 26617 18748
rect 26384 18708 26390 18720
rect 26605 18717 26617 18720
rect 26651 18717 26663 18751
rect 26605 18711 26663 18717
rect 26786 18708 26792 18760
rect 26844 18748 26850 18760
rect 26970 18748 26976 18760
rect 26844 18720 26976 18748
rect 26844 18708 26850 18720
rect 26970 18708 26976 18720
rect 27028 18708 27034 18760
rect 27065 18751 27123 18757
rect 27065 18717 27077 18751
rect 27111 18717 27123 18751
rect 27065 18711 27123 18717
rect 28077 18751 28135 18757
rect 28077 18717 28089 18751
rect 28123 18748 28135 18751
rect 29454 18748 29460 18760
rect 28123 18720 29460 18748
rect 28123 18717 28135 18720
rect 28077 18711 28135 18717
rect 26234 18680 26240 18692
rect 24872 18652 26240 18680
rect 26234 18640 26240 18652
rect 26292 18640 26298 18692
rect 27080 18680 27108 18711
rect 29454 18708 29460 18720
rect 29512 18708 29518 18760
rect 29730 18748 29736 18760
rect 29691 18720 29736 18748
rect 29730 18708 29736 18720
rect 29788 18708 29794 18760
rect 29914 18748 29920 18760
rect 29875 18720 29920 18748
rect 29914 18708 29920 18720
rect 29972 18708 29978 18760
rect 30190 18748 30196 18760
rect 30151 18720 30196 18748
rect 30190 18708 30196 18720
rect 30248 18708 30254 18760
rect 30834 18748 30840 18760
rect 30795 18720 30840 18748
rect 30834 18708 30840 18720
rect 30892 18708 30898 18760
rect 31018 18708 31024 18760
rect 31076 18748 31082 18760
rect 31113 18751 31171 18757
rect 31113 18748 31125 18751
rect 31076 18720 31125 18748
rect 31076 18708 31082 18720
rect 31113 18717 31125 18720
rect 31159 18717 31171 18751
rect 31113 18711 31171 18717
rect 31662 18708 31668 18760
rect 31720 18748 31726 18760
rect 31757 18751 31815 18757
rect 31757 18748 31769 18751
rect 31720 18720 31769 18748
rect 31720 18708 31726 18720
rect 31757 18717 31769 18720
rect 31803 18717 31815 18751
rect 31757 18711 31815 18717
rect 31846 18708 31852 18760
rect 31904 18748 31910 18760
rect 32674 18748 32680 18760
rect 31904 18720 31949 18748
rect 32635 18720 32680 18748
rect 31904 18708 31910 18720
rect 32674 18708 32680 18720
rect 32732 18708 32738 18760
rect 32858 18708 32864 18760
rect 32916 18748 32922 18760
rect 33045 18751 33103 18757
rect 33045 18748 33057 18751
rect 32916 18720 33057 18748
rect 32916 18708 32922 18720
rect 33045 18717 33057 18720
rect 33091 18717 33103 18751
rect 33045 18711 33103 18717
rect 33134 18708 33140 18760
rect 33192 18748 33198 18760
rect 33321 18751 33379 18757
rect 33192 18720 33237 18748
rect 33192 18708 33198 18720
rect 33321 18717 33333 18751
rect 33367 18748 33379 18751
rect 33781 18751 33839 18757
rect 33781 18748 33793 18751
rect 33367 18720 33793 18748
rect 33367 18717 33379 18720
rect 33321 18711 33379 18717
rect 33781 18717 33793 18720
rect 33827 18717 33839 18751
rect 33962 18748 33968 18760
rect 33923 18720 33968 18748
rect 33781 18711 33839 18717
rect 33962 18708 33968 18720
rect 34020 18708 34026 18760
rect 34790 18708 34796 18760
rect 34848 18748 34854 18760
rect 34885 18751 34943 18757
rect 34885 18748 34897 18751
rect 34848 18720 34897 18748
rect 34848 18708 34854 18720
rect 34885 18717 34897 18720
rect 34931 18717 34943 18751
rect 34885 18711 34943 18717
rect 30098 18689 30104 18692
rect 26804 18652 27108 18680
rect 29825 18683 29883 18689
rect 25130 18612 25136 18624
rect 24688 18584 25136 18612
rect 24397 18575 24455 18581
rect 25130 18572 25136 18584
rect 25188 18572 25194 18624
rect 26142 18572 26148 18624
rect 26200 18612 26206 18624
rect 26804 18612 26832 18652
rect 29825 18649 29837 18683
rect 29871 18649 29883 18683
rect 29825 18643 29883 18649
rect 30055 18683 30104 18689
rect 30055 18649 30067 18683
rect 30101 18649 30104 18683
rect 30055 18643 30104 18649
rect 26970 18612 26976 18624
rect 26200 18584 26832 18612
rect 26931 18584 26976 18612
rect 26200 18572 26206 18584
rect 26970 18572 26976 18584
rect 27028 18572 27034 18624
rect 28537 18615 28595 18621
rect 28537 18581 28549 18615
rect 28583 18612 28595 18615
rect 28718 18612 28724 18624
rect 28583 18584 28724 18612
rect 28583 18581 28595 18584
rect 28537 18575 28595 18581
rect 28718 18572 28724 18584
rect 28776 18572 28782 18624
rect 29840 18612 29868 18643
rect 30098 18640 30104 18643
rect 30156 18640 30162 18692
rect 33226 18680 33232 18692
rect 30576 18652 33232 18680
rect 30576 18612 30604 18652
rect 33226 18640 33232 18652
rect 33284 18640 33290 18692
rect 29840 18584 30604 18612
rect 31021 18615 31079 18621
rect 31021 18581 31033 18615
rect 31067 18612 31079 18615
rect 31110 18612 31116 18624
rect 31067 18584 31116 18612
rect 31067 18581 31079 18584
rect 31021 18575 31079 18581
rect 31110 18572 31116 18584
rect 31168 18572 31174 18624
rect 32125 18615 32183 18621
rect 32125 18581 32137 18615
rect 32171 18612 32183 18615
rect 32398 18612 32404 18624
rect 32171 18584 32404 18612
rect 32171 18581 32183 18584
rect 32125 18575 32183 18581
rect 32398 18572 32404 18584
rect 32456 18572 32462 18624
rect 32950 18572 32956 18624
rect 33008 18612 33014 18624
rect 33873 18615 33931 18621
rect 33873 18612 33885 18615
rect 33008 18584 33885 18612
rect 33008 18572 33014 18584
rect 33873 18581 33885 18584
rect 33919 18581 33931 18615
rect 33873 18575 33931 18581
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 12710 18408 12716 18420
rect 12671 18380 12716 18408
rect 12710 18368 12716 18380
rect 12768 18368 12774 18420
rect 13998 18408 14004 18420
rect 13372 18380 14004 18408
rect 9668 18343 9726 18349
rect 9668 18309 9680 18343
rect 9714 18340 9726 18343
rect 10502 18340 10508 18352
rect 9714 18312 10508 18340
rect 9714 18309 9726 18312
rect 9668 18303 9726 18309
rect 10502 18300 10508 18312
rect 10560 18300 10566 18352
rect 11977 18343 12035 18349
rect 11977 18309 11989 18343
rect 12023 18309 12035 18343
rect 11977 18303 12035 18309
rect 12161 18343 12219 18349
rect 12161 18309 12173 18343
rect 12207 18340 12219 18343
rect 12434 18340 12440 18352
rect 12207 18312 12440 18340
rect 12207 18309 12219 18312
rect 12161 18303 12219 18309
rect 9398 18272 9404 18284
rect 9311 18244 9404 18272
rect 9398 18232 9404 18244
rect 9456 18272 9462 18284
rect 11882 18272 11888 18284
rect 9456 18244 11888 18272
rect 9456 18232 9462 18244
rect 11882 18232 11888 18244
rect 11940 18232 11946 18284
rect 10778 18136 10784 18148
rect 10691 18108 10784 18136
rect 10778 18096 10784 18108
rect 10836 18136 10842 18148
rect 11992 18136 12020 18303
rect 12434 18300 12440 18312
rect 12492 18300 12498 18352
rect 12897 18275 12955 18281
rect 12897 18241 12909 18275
rect 12943 18272 12955 18275
rect 12986 18272 12992 18284
rect 12943 18244 12992 18272
rect 12943 18241 12955 18244
rect 12897 18235 12955 18241
rect 12986 18232 12992 18244
rect 13044 18232 13050 18284
rect 13170 18272 13176 18284
rect 13131 18244 13176 18272
rect 13170 18232 13176 18244
rect 13228 18232 13234 18284
rect 13372 18281 13400 18380
rect 13998 18368 14004 18380
rect 14056 18368 14062 18420
rect 16117 18411 16175 18417
rect 16117 18377 16129 18411
rect 16163 18408 16175 18411
rect 16574 18408 16580 18420
rect 16163 18380 16580 18408
rect 16163 18377 16175 18380
rect 16117 18371 16175 18377
rect 16574 18368 16580 18380
rect 16632 18368 16638 18420
rect 16942 18368 16948 18420
rect 17000 18408 17006 18420
rect 18049 18411 18107 18417
rect 18049 18408 18061 18411
rect 17000 18380 18061 18408
rect 17000 18368 17006 18380
rect 18049 18377 18061 18380
rect 18095 18377 18107 18411
rect 18049 18371 18107 18377
rect 18138 18368 18144 18420
rect 18196 18408 18202 18420
rect 20993 18411 21051 18417
rect 20993 18408 21005 18411
rect 18196 18380 21005 18408
rect 18196 18368 18202 18380
rect 20993 18377 21005 18380
rect 21039 18377 21051 18411
rect 20993 18371 21051 18377
rect 23658 18368 23664 18420
rect 23716 18408 23722 18420
rect 23753 18411 23811 18417
rect 23753 18408 23765 18411
rect 23716 18380 23765 18408
rect 23716 18368 23722 18380
rect 23753 18377 23765 18380
rect 23799 18377 23811 18411
rect 25590 18408 25596 18420
rect 25551 18380 25596 18408
rect 23753 18371 23811 18377
rect 25590 18368 25596 18380
rect 25648 18368 25654 18420
rect 25866 18368 25872 18420
rect 25924 18408 25930 18420
rect 26237 18411 26295 18417
rect 26237 18408 26249 18411
rect 25924 18380 26249 18408
rect 25924 18368 25930 18380
rect 26237 18377 26249 18380
rect 26283 18377 26295 18411
rect 26237 18371 26295 18377
rect 26970 18368 26976 18420
rect 27028 18408 27034 18420
rect 29181 18411 29239 18417
rect 29181 18408 29193 18411
rect 27028 18380 29193 18408
rect 27028 18368 27034 18380
rect 29181 18377 29193 18380
rect 29227 18377 29239 18411
rect 29181 18371 29239 18377
rect 29730 18368 29736 18420
rect 29788 18408 29794 18420
rect 31202 18408 31208 18420
rect 29788 18380 31208 18408
rect 29788 18368 29794 18380
rect 31202 18368 31208 18380
rect 31260 18368 31266 18420
rect 32493 18411 32551 18417
rect 32493 18377 32505 18411
rect 32539 18408 32551 18411
rect 32674 18408 32680 18420
rect 32539 18380 32680 18408
rect 32539 18377 32551 18380
rect 32493 18371 32551 18377
rect 32674 18368 32680 18380
rect 32732 18368 32738 18420
rect 33226 18368 33232 18420
rect 33284 18408 33290 18420
rect 33321 18411 33379 18417
rect 33321 18408 33333 18411
rect 33284 18380 33333 18408
rect 33284 18368 33290 18380
rect 33321 18377 33333 18380
rect 33367 18377 33379 18411
rect 33321 18371 33379 18377
rect 13814 18300 13820 18352
rect 13872 18340 13878 18352
rect 13909 18343 13967 18349
rect 13909 18340 13921 18343
rect 13872 18312 13921 18340
rect 13872 18300 13878 18312
rect 13909 18309 13921 18312
rect 13955 18309 13967 18343
rect 15930 18340 15936 18352
rect 15891 18312 15936 18340
rect 13909 18303 13967 18309
rect 15930 18300 15936 18312
rect 15988 18300 15994 18352
rect 17034 18340 17040 18352
rect 16995 18312 17040 18340
rect 17034 18300 17040 18312
rect 17092 18300 17098 18352
rect 17126 18300 17132 18352
rect 17184 18340 17190 18352
rect 17957 18343 18015 18349
rect 17184 18312 17229 18340
rect 17184 18300 17190 18312
rect 17957 18309 17969 18343
rect 18003 18340 18015 18343
rect 19334 18340 19340 18352
rect 18003 18312 19340 18340
rect 18003 18309 18015 18312
rect 17957 18303 18015 18309
rect 19334 18300 19340 18312
rect 19392 18300 19398 18352
rect 23474 18340 23480 18352
rect 20456 18312 23480 18340
rect 13357 18275 13415 18281
rect 13357 18241 13369 18275
rect 13403 18241 13415 18275
rect 13357 18235 13415 18241
rect 15105 18275 15163 18281
rect 15105 18241 15117 18275
rect 15151 18241 15163 18275
rect 15286 18272 15292 18284
rect 15247 18244 15292 18272
rect 15105 18235 15163 18241
rect 10836 18108 12020 18136
rect 10836 18096 10842 18108
rect 15120 18068 15148 18235
rect 15286 18232 15292 18244
rect 15344 18232 15350 18284
rect 15749 18275 15807 18281
rect 15749 18241 15761 18275
rect 15795 18272 15807 18275
rect 16482 18272 16488 18284
rect 15795 18244 16488 18272
rect 15795 18241 15807 18244
rect 15749 18235 15807 18241
rect 16482 18232 16488 18244
rect 16540 18232 16546 18284
rect 16853 18275 16911 18281
rect 16853 18241 16865 18275
rect 16899 18241 16911 18275
rect 16853 18235 16911 18241
rect 17221 18275 17279 18281
rect 17221 18241 17233 18275
rect 17267 18241 17279 18275
rect 17221 18235 17279 18241
rect 15197 18207 15255 18213
rect 15197 18173 15209 18207
rect 15243 18204 15255 18207
rect 16390 18204 16396 18216
rect 15243 18176 16396 18204
rect 15243 18173 15255 18176
rect 15197 18167 15255 18173
rect 16390 18164 16396 18176
rect 16448 18204 16454 18216
rect 16868 18204 16896 18235
rect 16448 18176 16896 18204
rect 16448 18164 16454 18176
rect 17034 18164 17040 18216
rect 17092 18204 17098 18216
rect 17236 18204 17264 18235
rect 18230 18232 18236 18284
rect 18288 18272 18294 18284
rect 18693 18275 18751 18281
rect 18693 18272 18705 18275
rect 18288 18244 18705 18272
rect 18288 18232 18294 18244
rect 18693 18241 18705 18244
rect 18739 18241 18751 18275
rect 18693 18235 18751 18241
rect 18969 18275 19027 18281
rect 18969 18241 18981 18275
rect 19015 18272 19027 18275
rect 19242 18272 19248 18284
rect 19015 18244 19248 18272
rect 19015 18241 19027 18244
rect 18969 18235 19027 18241
rect 19242 18232 19248 18244
rect 19300 18232 19306 18284
rect 19981 18275 20039 18281
rect 19981 18241 19993 18275
rect 20027 18272 20039 18275
rect 20162 18272 20168 18284
rect 20027 18244 20168 18272
rect 20027 18241 20039 18244
rect 19981 18235 20039 18241
rect 20162 18232 20168 18244
rect 20220 18232 20226 18284
rect 20255 18275 20313 18281
rect 20255 18241 20267 18275
rect 20301 18270 20313 18275
rect 20456 18270 20484 18312
rect 23474 18300 23480 18312
rect 23532 18300 23538 18352
rect 25958 18340 25964 18352
rect 25516 18312 25964 18340
rect 21818 18272 21824 18284
rect 20301 18242 20484 18270
rect 21779 18244 21824 18272
rect 20301 18241 20313 18242
rect 20255 18235 20313 18241
rect 21818 18232 21824 18244
rect 21876 18232 21882 18284
rect 22002 18272 22008 18284
rect 21963 18244 22008 18272
rect 22002 18232 22008 18244
rect 22060 18232 22066 18284
rect 23017 18275 23075 18281
rect 23017 18241 23029 18275
rect 23063 18272 23075 18275
rect 23566 18272 23572 18284
rect 23063 18244 23572 18272
rect 23063 18241 23075 18244
rect 23017 18235 23075 18241
rect 23566 18232 23572 18244
rect 23624 18232 23630 18284
rect 24397 18275 24455 18281
rect 24397 18241 24409 18275
rect 24443 18272 24455 18275
rect 24762 18272 24768 18284
rect 24443 18244 24768 18272
rect 24443 18241 24455 18244
rect 24397 18235 24455 18241
rect 24762 18232 24768 18244
rect 24820 18232 24826 18284
rect 25516 18281 25544 18312
rect 25958 18300 25964 18312
rect 26016 18300 26022 18352
rect 26329 18343 26387 18349
rect 26329 18309 26341 18343
rect 26375 18340 26387 18343
rect 26786 18340 26792 18352
rect 26375 18312 26792 18340
rect 26375 18309 26387 18312
rect 26329 18303 26387 18309
rect 26786 18300 26792 18312
rect 26844 18300 26850 18352
rect 25501 18275 25559 18281
rect 25501 18241 25513 18275
rect 25547 18241 25559 18275
rect 25501 18235 25559 18241
rect 25685 18275 25743 18281
rect 25685 18241 25697 18275
rect 25731 18272 25743 18275
rect 25774 18272 25780 18284
rect 25731 18244 25780 18272
rect 25731 18241 25743 18244
rect 25685 18235 25743 18241
rect 25774 18232 25780 18244
rect 25832 18232 25838 18284
rect 26142 18272 26148 18284
rect 26055 18244 26148 18272
rect 26142 18232 26148 18244
rect 26200 18232 26206 18284
rect 26421 18275 26479 18281
rect 26421 18241 26433 18275
rect 26467 18272 26479 18275
rect 26988 18272 27016 18368
rect 30190 18340 30196 18352
rect 26467 18244 27016 18272
rect 27080 18312 30196 18340
rect 26467 18241 26479 18244
rect 26421 18235 26479 18241
rect 22738 18204 22744 18216
rect 17092 18176 17264 18204
rect 22699 18176 22744 18204
rect 17092 18164 17098 18176
rect 22738 18164 22744 18176
rect 22796 18164 22802 18216
rect 25314 18164 25320 18216
rect 25372 18204 25378 18216
rect 26160 18204 26188 18232
rect 25372 18176 26188 18204
rect 25372 18164 25378 18176
rect 16758 18096 16764 18148
rect 16816 18136 16822 18148
rect 17052 18136 17080 18164
rect 16816 18108 17080 18136
rect 16816 18096 16822 18108
rect 17218 18096 17224 18148
rect 17276 18136 17282 18148
rect 17405 18139 17463 18145
rect 17405 18136 17417 18139
rect 17276 18108 17417 18136
rect 17276 18096 17282 18108
rect 17405 18105 17417 18108
rect 17451 18105 17463 18139
rect 17405 18099 17463 18105
rect 26050 18096 26056 18148
rect 26108 18136 26114 18148
rect 27080 18136 27108 18312
rect 30190 18300 30196 18312
rect 30248 18300 30254 18352
rect 31386 18340 31392 18352
rect 30760 18312 31392 18340
rect 27893 18275 27951 18281
rect 27893 18241 27905 18275
rect 27939 18241 27951 18275
rect 28718 18272 28724 18284
rect 27893 18235 27951 18241
rect 28000 18244 28724 18272
rect 26108 18108 27108 18136
rect 27908 18136 27936 18235
rect 28000 18213 28028 18244
rect 28718 18232 28724 18244
rect 28776 18232 28782 18284
rect 30760 18213 30788 18312
rect 31386 18300 31392 18312
rect 31444 18300 31450 18352
rect 32398 18300 32404 18352
rect 32456 18340 32462 18352
rect 33137 18343 33195 18349
rect 33137 18340 33149 18343
rect 32456 18312 33149 18340
rect 32456 18300 32462 18312
rect 33137 18309 33149 18312
rect 33183 18309 33195 18343
rect 33137 18303 33195 18309
rect 30837 18275 30895 18281
rect 30837 18241 30849 18275
rect 30883 18272 30895 18275
rect 31294 18272 31300 18284
rect 30883 18244 31300 18272
rect 30883 18241 30895 18244
rect 30837 18235 30895 18241
rect 31294 18232 31300 18244
rect 31352 18232 31358 18284
rect 31662 18232 31668 18284
rect 31720 18272 31726 18284
rect 32122 18272 32128 18284
rect 31720 18244 32128 18272
rect 31720 18232 31726 18244
rect 32122 18232 32128 18244
rect 32180 18232 32186 18284
rect 32950 18272 32956 18284
rect 32911 18244 32956 18272
rect 32950 18232 32956 18244
rect 33008 18232 33014 18284
rect 33336 18272 33364 18371
rect 33962 18368 33968 18420
rect 34020 18368 34026 18420
rect 34974 18408 34980 18420
rect 34935 18380 34980 18408
rect 34974 18368 34980 18380
rect 35032 18368 35038 18420
rect 33980 18340 34008 18368
rect 33980 18312 34836 18340
rect 33965 18275 34023 18281
rect 33965 18272 33977 18275
rect 33336 18244 33977 18272
rect 33965 18241 33977 18244
rect 34011 18272 34023 18275
rect 34146 18272 34152 18284
rect 34011 18244 34152 18272
rect 34011 18241 34023 18244
rect 33965 18235 34023 18241
rect 34146 18232 34152 18244
rect 34204 18232 34210 18284
rect 34808 18281 34836 18312
rect 34793 18275 34851 18281
rect 34793 18241 34805 18275
rect 34839 18241 34851 18275
rect 34793 18235 34851 18241
rect 34977 18275 35035 18281
rect 34977 18241 34989 18275
rect 35023 18272 35035 18275
rect 35342 18272 35348 18284
rect 35023 18244 35348 18272
rect 35023 18241 35035 18244
rect 34977 18235 35035 18241
rect 35342 18232 35348 18244
rect 35400 18232 35406 18284
rect 27985 18207 28043 18213
rect 27985 18173 27997 18207
rect 28031 18173 28043 18207
rect 27985 18167 28043 18173
rect 30745 18207 30803 18213
rect 30745 18173 30757 18207
rect 30791 18173 30803 18207
rect 30745 18167 30803 18173
rect 31110 18164 31116 18216
rect 31168 18204 31174 18216
rect 31478 18204 31484 18216
rect 31168 18176 31484 18204
rect 31168 18164 31174 18176
rect 31478 18164 31484 18176
rect 31536 18204 31542 18216
rect 32217 18207 32275 18213
rect 32217 18204 32229 18207
rect 31536 18176 32229 18204
rect 31536 18164 31542 18176
rect 32217 18173 32229 18176
rect 32263 18173 32275 18207
rect 34054 18204 34060 18216
rect 34015 18176 34060 18204
rect 32217 18167 32275 18173
rect 34054 18164 34060 18176
rect 34112 18164 34118 18216
rect 34330 18204 34336 18216
rect 34291 18176 34336 18204
rect 34330 18164 34336 18176
rect 34388 18164 34394 18216
rect 27908 18108 28304 18136
rect 26108 18096 26114 18108
rect 18230 18068 18236 18080
rect 15120 18040 18236 18068
rect 18230 18028 18236 18040
rect 18288 18028 18294 18080
rect 19150 18028 19156 18080
rect 19208 18068 19214 18080
rect 21821 18071 21879 18077
rect 21821 18068 21833 18071
rect 19208 18040 21833 18068
rect 19208 18028 19214 18040
rect 21821 18037 21833 18040
rect 21867 18037 21879 18071
rect 21821 18031 21879 18037
rect 24213 18071 24271 18077
rect 24213 18037 24225 18071
rect 24259 18068 24271 18071
rect 25222 18068 25228 18080
rect 24259 18040 25228 18068
rect 24259 18037 24271 18040
rect 24213 18031 24271 18037
rect 25222 18028 25228 18040
rect 25280 18028 25286 18080
rect 27982 18028 27988 18080
rect 28040 18068 28046 18080
rect 28169 18071 28227 18077
rect 28169 18068 28181 18071
rect 28040 18040 28181 18068
rect 28040 18028 28046 18040
rect 28169 18037 28181 18040
rect 28215 18037 28227 18071
rect 28276 18068 28304 18108
rect 28626 18096 28632 18148
rect 28684 18136 28690 18148
rect 31205 18139 31263 18145
rect 31205 18136 31217 18139
rect 28684 18108 31217 18136
rect 28684 18096 28690 18108
rect 31205 18105 31217 18108
rect 31251 18105 31263 18139
rect 31205 18099 31263 18105
rect 28905 18071 28963 18077
rect 28905 18068 28917 18071
rect 28276 18040 28917 18068
rect 28169 18031 28227 18037
rect 28905 18037 28917 18040
rect 28951 18068 28963 18071
rect 29178 18068 29184 18080
rect 28951 18040 29184 18068
rect 28951 18037 28963 18040
rect 28905 18031 28963 18037
rect 29178 18028 29184 18040
rect 29236 18028 29242 18080
rect 31754 18028 31760 18080
rect 31812 18068 31818 18080
rect 32125 18071 32183 18077
rect 32125 18068 32137 18071
rect 31812 18040 32137 18068
rect 31812 18028 31818 18040
rect 32125 18037 32137 18040
rect 32171 18037 32183 18071
rect 32125 18031 32183 18037
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 10594 17864 10600 17876
rect 10555 17836 10600 17864
rect 10594 17824 10600 17836
rect 10652 17824 10658 17876
rect 11054 17824 11060 17876
rect 11112 17864 11118 17876
rect 11333 17867 11391 17873
rect 11333 17864 11345 17867
rect 11112 17836 11345 17864
rect 11112 17824 11118 17836
rect 11333 17833 11345 17836
rect 11379 17833 11391 17867
rect 14274 17864 14280 17876
rect 14235 17836 14280 17864
rect 11333 17827 11391 17833
rect 14274 17824 14280 17836
rect 14332 17824 14338 17876
rect 20162 17824 20168 17876
rect 20220 17864 20226 17876
rect 21818 17864 21824 17876
rect 20220 17836 21824 17864
rect 20220 17824 20226 17836
rect 18601 17799 18659 17805
rect 18601 17796 18613 17799
rect 15396 17768 18613 17796
rect 15396 17737 15424 17768
rect 18601 17765 18613 17768
rect 18647 17796 18659 17799
rect 18690 17796 18696 17808
rect 18647 17768 18696 17796
rect 18647 17765 18659 17768
rect 18601 17759 18659 17765
rect 18690 17756 18696 17768
rect 18748 17756 18754 17808
rect 21008 17805 21036 17836
rect 21818 17824 21824 17836
rect 21876 17824 21882 17876
rect 21910 17824 21916 17876
rect 21968 17864 21974 17876
rect 24578 17864 24584 17876
rect 21968 17836 23704 17864
rect 24539 17836 24584 17864
rect 21968 17824 21974 17836
rect 20257 17799 20315 17805
rect 20257 17765 20269 17799
rect 20303 17765 20315 17799
rect 20257 17759 20315 17765
rect 20993 17799 21051 17805
rect 20993 17765 21005 17799
rect 21039 17765 21051 17799
rect 20993 17759 21051 17765
rect 23569 17799 23627 17805
rect 23569 17765 23581 17799
rect 23615 17765 23627 17799
rect 23569 17759 23627 17765
rect 15381 17731 15439 17737
rect 15381 17697 15393 17731
rect 15427 17697 15439 17731
rect 15381 17691 15439 17697
rect 15565 17731 15623 17737
rect 15565 17697 15577 17731
rect 15611 17728 15623 17731
rect 15838 17728 15844 17740
rect 15611 17700 15844 17728
rect 15611 17697 15623 17700
rect 15565 17691 15623 17697
rect 15838 17688 15844 17700
rect 15896 17688 15902 17740
rect 16206 17728 16212 17740
rect 16167 17700 16212 17728
rect 16206 17688 16212 17700
rect 16264 17688 16270 17740
rect 16485 17731 16543 17737
rect 16485 17697 16497 17731
rect 16531 17728 16543 17731
rect 17497 17731 17555 17737
rect 17497 17728 17509 17731
rect 16531 17700 17509 17728
rect 16531 17697 16543 17700
rect 16485 17691 16543 17697
rect 17497 17697 17509 17700
rect 17543 17728 17555 17731
rect 20272 17728 20300 17759
rect 23584 17728 23612 17759
rect 17543 17700 18092 17728
rect 20272 17700 20944 17728
rect 17543 17697 17555 17700
rect 17497 17691 17555 17697
rect 18064 17672 18092 17700
rect 9766 17620 9772 17672
rect 9824 17660 9830 17672
rect 10594 17660 10600 17672
rect 9824 17632 10600 17660
rect 9824 17620 9830 17632
rect 10594 17620 10600 17632
rect 10652 17620 10658 17672
rect 10778 17660 10784 17672
rect 10739 17632 10784 17660
rect 10778 17620 10784 17632
rect 10836 17620 10842 17672
rect 11238 17660 11244 17672
rect 11199 17632 11244 17660
rect 11238 17620 11244 17632
rect 11296 17620 11302 17672
rect 11425 17663 11483 17669
rect 11425 17629 11437 17663
rect 11471 17660 11483 17663
rect 12158 17660 12164 17672
rect 11471 17632 12164 17660
rect 11471 17629 11483 17632
rect 11425 17623 11483 17629
rect 12158 17620 12164 17632
rect 12216 17620 12222 17672
rect 14461 17663 14519 17669
rect 14461 17629 14473 17663
rect 14507 17660 14519 17663
rect 15010 17660 15016 17672
rect 14507 17632 15016 17660
rect 14507 17629 14519 17632
rect 14461 17623 14519 17629
rect 15010 17620 15016 17632
rect 15068 17620 15074 17672
rect 17681 17663 17739 17669
rect 17681 17629 17693 17663
rect 17727 17629 17739 17663
rect 17681 17623 17739 17629
rect 15289 17595 15347 17601
rect 15289 17561 15301 17595
rect 15335 17592 15347 17595
rect 16942 17592 16948 17604
rect 15335 17564 16948 17592
rect 15335 17561 15347 17564
rect 15289 17555 15347 17561
rect 16942 17552 16948 17564
rect 17000 17552 17006 17604
rect 17696 17592 17724 17623
rect 18046 17620 18052 17672
rect 18104 17660 18110 17672
rect 18417 17663 18475 17669
rect 18417 17660 18429 17663
rect 18104 17632 18429 17660
rect 18104 17620 18110 17632
rect 18417 17629 18429 17632
rect 18463 17629 18475 17663
rect 18417 17623 18475 17629
rect 19245 17663 19303 17669
rect 19245 17629 19257 17663
rect 19291 17629 19303 17663
rect 19518 17660 19524 17672
rect 19479 17632 19524 17660
rect 19245 17623 19303 17629
rect 18322 17592 18328 17604
rect 17696 17564 18328 17592
rect 18322 17552 18328 17564
rect 18380 17592 18386 17604
rect 19260 17592 19288 17623
rect 19518 17620 19524 17632
rect 19576 17620 19582 17672
rect 20806 17660 20812 17672
rect 20767 17632 20812 17660
rect 20806 17620 20812 17632
rect 20864 17620 20870 17672
rect 20916 17669 20944 17700
rect 22848 17700 23612 17728
rect 23676 17728 23704 17836
rect 24578 17824 24584 17836
rect 24636 17824 24642 17876
rect 24762 17864 24768 17876
rect 24723 17836 24768 17864
rect 24762 17824 24768 17836
rect 24820 17824 24826 17876
rect 27709 17867 27767 17873
rect 27709 17833 27721 17867
rect 27755 17864 27767 17867
rect 30098 17864 30104 17876
rect 27755 17836 30104 17864
rect 27755 17833 27767 17836
rect 27709 17827 27767 17833
rect 30098 17824 30104 17836
rect 30156 17824 30162 17876
rect 30374 17824 30380 17876
rect 30432 17864 30438 17876
rect 30653 17867 30711 17873
rect 30653 17864 30665 17867
rect 30432 17836 30665 17864
rect 30432 17824 30438 17836
rect 30653 17833 30665 17836
rect 30699 17833 30711 17867
rect 31386 17864 31392 17876
rect 31347 17836 31392 17864
rect 30653 17827 30711 17833
rect 23750 17756 23756 17808
rect 23808 17796 23814 17808
rect 25869 17799 25927 17805
rect 25869 17796 25881 17799
rect 23808 17768 25881 17796
rect 23808 17756 23814 17768
rect 25869 17765 25881 17768
rect 25915 17765 25927 17799
rect 25869 17759 25927 17765
rect 26786 17756 26792 17808
rect 26844 17796 26850 17808
rect 26844 17768 27384 17796
rect 26844 17756 26850 17768
rect 27246 17728 27252 17740
rect 23676 17700 24440 17728
rect 27207 17700 27252 17728
rect 20901 17663 20959 17669
rect 20901 17629 20913 17663
rect 20947 17629 20959 17663
rect 20901 17623 20959 17629
rect 21450 17620 21456 17672
rect 21508 17660 21514 17672
rect 21545 17663 21603 17669
rect 21545 17660 21557 17663
rect 21508 17632 21557 17660
rect 21508 17620 21514 17632
rect 21545 17629 21557 17632
rect 21591 17629 21603 17663
rect 21545 17623 21603 17629
rect 21821 17663 21879 17669
rect 21821 17629 21833 17663
rect 21867 17660 21879 17663
rect 22848 17660 22876 17700
rect 21867 17632 22876 17660
rect 23017 17663 23075 17669
rect 21867 17629 21879 17632
rect 21821 17623 21879 17629
rect 23017 17629 23029 17663
rect 23063 17629 23075 17663
rect 23290 17660 23296 17672
rect 23251 17632 23296 17660
rect 23017 17623 23075 17629
rect 18380 17564 19288 17592
rect 18380 17552 18386 17564
rect 19334 17552 19340 17604
rect 19392 17592 19398 17604
rect 19536 17592 19564 17620
rect 19392 17564 19564 17592
rect 19392 17552 19398 17564
rect 20438 17552 20444 17604
rect 20496 17592 20502 17604
rect 23032 17592 23060 17623
rect 23290 17620 23296 17632
rect 23348 17620 23354 17672
rect 23382 17620 23388 17672
rect 23440 17660 23446 17672
rect 23440 17632 23485 17660
rect 23440 17620 23446 17632
rect 24412 17601 24440 17700
rect 27246 17688 27252 17700
rect 27304 17688 27310 17740
rect 24670 17620 24676 17672
rect 24728 17660 24734 17672
rect 25498 17660 25504 17672
rect 24728 17632 25504 17660
rect 24728 17620 24734 17632
rect 25498 17620 25504 17632
rect 25556 17660 25562 17672
rect 25869 17663 25927 17669
rect 25869 17660 25881 17663
rect 25556 17632 25881 17660
rect 25556 17620 25562 17632
rect 25869 17629 25881 17632
rect 25915 17629 25927 17663
rect 25869 17623 25927 17629
rect 26145 17663 26203 17669
rect 26145 17629 26157 17663
rect 26191 17660 26203 17663
rect 27154 17660 27160 17672
rect 26191 17632 27160 17660
rect 26191 17629 26203 17632
rect 26145 17623 26203 17629
rect 27154 17620 27160 17632
rect 27212 17620 27218 17672
rect 27356 17669 27384 17768
rect 30668 17728 30696 17827
rect 31386 17824 31392 17836
rect 31444 17824 31450 17876
rect 31202 17756 31208 17808
rect 31260 17796 31266 17808
rect 32309 17799 32367 17805
rect 32309 17796 32321 17799
rect 31260 17768 32321 17796
rect 31260 17756 31266 17768
rect 32309 17765 32321 17768
rect 32355 17765 32367 17799
rect 32309 17759 32367 17765
rect 32950 17728 32956 17740
rect 30668 17700 31754 17728
rect 27341 17663 27399 17669
rect 27341 17629 27353 17663
rect 27387 17629 27399 17663
rect 27341 17623 27399 17629
rect 30561 17663 30619 17669
rect 30561 17629 30573 17663
rect 30607 17629 30619 17663
rect 30834 17660 30840 17672
rect 30795 17632 30840 17660
rect 30561 17623 30619 17629
rect 20496 17564 23060 17592
rect 23201 17595 23259 17601
rect 20496 17552 20502 17564
rect 23201 17561 23213 17595
rect 23247 17561 23259 17595
rect 23201 17555 23259 17561
rect 24397 17595 24455 17601
rect 24397 17561 24409 17595
rect 24443 17561 24455 17595
rect 26418 17592 26424 17604
rect 24397 17555 24455 17561
rect 25976 17564 26424 17592
rect 14918 17524 14924 17536
rect 14879 17496 14924 17524
rect 14918 17484 14924 17496
rect 14976 17484 14982 17536
rect 17862 17524 17868 17536
rect 17823 17496 17868 17524
rect 17862 17484 17868 17496
rect 17920 17484 17926 17536
rect 19058 17484 19064 17536
rect 19116 17524 19122 17536
rect 20162 17524 20168 17536
rect 19116 17496 20168 17524
rect 19116 17484 19122 17496
rect 20162 17484 20168 17496
rect 20220 17484 20226 17536
rect 22554 17524 22560 17536
rect 22515 17496 22560 17524
rect 22554 17484 22560 17496
rect 22612 17484 22618 17536
rect 22646 17484 22652 17536
rect 22704 17524 22710 17536
rect 23216 17524 23244 17555
rect 22704 17496 23244 17524
rect 24607 17527 24665 17533
rect 22704 17484 22710 17496
rect 24607 17493 24619 17527
rect 24653 17524 24665 17527
rect 25976 17524 26004 17564
rect 26418 17552 26424 17564
rect 26476 17552 26482 17604
rect 24653 17496 26004 17524
rect 26053 17527 26111 17533
rect 24653 17493 24665 17496
rect 24607 17487 24665 17493
rect 26053 17493 26065 17527
rect 26099 17524 26111 17527
rect 27798 17524 27804 17536
rect 26099 17496 27804 17524
rect 26099 17493 26111 17496
rect 26053 17487 26111 17493
rect 27798 17484 27804 17496
rect 27856 17484 27862 17536
rect 30576 17524 30604 17623
rect 30834 17620 30840 17632
rect 30892 17620 30898 17672
rect 31312 17669 31340 17700
rect 31297 17663 31355 17669
rect 31297 17629 31309 17663
rect 31343 17629 31355 17663
rect 31478 17660 31484 17672
rect 31439 17632 31484 17660
rect 31297 17623 31355 17629
rect 31478 17620 31484 17632
rect 31536 17620 31542 17672
rect 30745 17595 30803 17601
rect 30745 17561 30757 17595
rect 30791 17592 30803 17595
rect 31496 17592 31524 17620
rect 30791 17564 31524 17592
rect 31726 17592 31754 17700
rect 32232 17700 32956 17728
rect 32232 17669 32260 17700
rect 32950 17688 32956 17700
rect 33008 17688 33014 17740
rect 32217 17663 32275 17669
rect 32217 17629 32229 17663
rect 32263 17629 32275 17663
rect 32398 17660 32404 17672
rect 32359 17632 32404 17660
rect 32217 17623 32275 17629
rect 32398 17620 32404 17632
rect 32456 17620 32462 17672
rect 31846 17592 31852 17604
rect 31726 17564 31852 17592
rect 30791 17561 30803 17564
rect 30745 17555 30803 17561
rect 31846 17552 31852 17564
rect 31904 17552 31910 17604
rect 31018 17524 31024 17536
rect 30576 17496 31024 17524
rect 31018 17484 31024 17496
rect 31076 17484 31082 17536
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 12342 17320 12348 17332
rect 12303 17292 12348 17320
rect 12342 17280 12348 17292
rect 12400 17280 12406 17332
rect 15565 17323 15623 17329
rect 15565 17289 15577 17323
rect 15611 17320 15623 17323
rect 16206 17320 16212 17332
rect 15611 17292 16212 17320
rect 15611 17289 15623 17292
rect 15565 17283 15623 17289
rect 16206 17280 16212 17292
rect 16264 17280 16270 17332
rect 21177 17323 21235 17329
rect 21177 17320 21189 17323
rect 16684 17292 21189 17320
rect 10413 17255 10471 17261
rect 10413 17221 10425 17255
rect 10459 17252 10471 17255
rect 11330 17252 11336 17264
rect 10459 17224 11336 17252
rect 10459 17221 10471 17224
rect 10413 17215 10471 17221
rect 11330 17212 11336 17224
rect 11388 17212 11394 17264
rect 12802 17252 12808 17264
rect 12544 17224 12808 17252
rect 10229 17187 10287 17193
rect 10229 17153 10241 17187
rect 10275 17184 10287 17187
rect 10318 17184 10324 17196
rect 10275 17156 10324 17184
rect 10275 17153 10287 17156
rect 10229 17147 10287 17153
rect 10318 17144 10324 17156
rect 10376 17144 10382 17196
rect 12544 17193 12572 17224
rect 12802 17212 12808 17224
rect 12860 17252 12866 17264
rect 13725 17255 13783 17261
rect 13725 17252 13737 17255
rect 12860 17224 13737 17252
rect 12860 17212 12866 17224
rect 13725 17221 13737 17224
rect 13771 17221 13783 17255
rect 13725 17215 13783 17221
rect 14182 17212 14188 17264
rect 14240 17252 14246 17264
rect 14240 17224 15240 17252
rect 14240 17212 14246 17224
rect 12529 17187 12587 17193
rect 12529 17153 12541 17187
rect 12575 17153 12587 17187
rect 12529 17147 12587 17153
rect 12621 17187 12679 17193
rect 12621 17153 12633 17187
rect 12667 17184 12679 17187
rect 12710 17184 12716 17196
rect 12667 17156 12716 17184
rect 12667 17153 12679 17156
rect 12621 17147 12679 17153
rect 12710 17144 12716 17156
rect 12768 17144 12774 17196
rect 12894 17184 12900 17196
rect 12855 17156 12900 17184
rect 12894 17144 12900 17156
rect 12952 17144 12958 17196
rect 13541 17187 13599 17193
rect 13541 17153 13553 17187
rect 13587 17184 13599 17187
rect 14090 17184 14096 17196
rect 13587 17156 14096 17184
rect 13587 17153 13599 17156
rect 13541 17147 13599 17153
rect 14090 17144 14096 17156
rect 14148 17144 14154 17196
rect 14452 17187 14510 17193
rect 14452 17153 14464 17187
rect 14498 17184 14510 17187
rect 14734 17184 14740 17196
rect 14498 17156 14740 17184
rect 14498 17153 14510 17156
rect 14452 17147 14510 17153
rect 14734 17144 14740 17156
rect 14792 17144 14798 17196
rect 13078 17076 13084 17128
rect 13136 17116 13142 17128
rect 13357 17119 13415 17125
rect 13357 17116 13369 17119
rect 13136 17088 13369 17116
rect 13136 17076 13142 17088
rect 13357 17085 13369 17088
rect 13403 17085 13415 17119
rect 14182 17116 14188 17128
rect 14143 17088 14188 17116
rect 13357 17079 13415 17085
rect 14182 17076 14188 17088
rect 14240 17076 14246 17128
rect 15212 17116 15240 17224
rect 16684 17193 16712 17292
rect 21177 17289 21189 17292
rect 21223 17289 21235 17323
rect 25961 17323 26019 17329
rect 25961 17320 25973 17323
rect 21177 17283 21235 17289
rect 22066 17292 25973 17320
rect 16850 17252 16856 17264
rect 16811 17224 16856 17252
rect 16850 17212 16856 17224
rect 16908 17212 16914 17264
rect 16942 17212 16948 17264
rect 17000 17252 17006 17264
rect 17000 17224 17045 17252
rect 17000 17212 17006 17224
rect 17126 17212 17132 17264
rect 17184 17252 17190 17264
rect 17681 17255 17739 17261
rect 17681 17252 17693 17255
rect 17184 17224 17693 17252
rect 17184 17212 17190 17224
rect 17681 17221 17693 17224
rect 17727 17221 17739 17255
rect 17681 17215 17739 17221
rect 17897 17255 17955 17261
rect 17897 17221 17909 17255
rect 17943 17252 17955 17255
rect 18322 17252 18328 17264
rect 17943 17224 18328 17252
rect 17943 17221 17955 17224
rect 17897 17215 17955 17221
rect 18322 17212 18328 17224
rect 18380 17212 18386 17264
rect 20257 17255 20315 17261
rect 20257 17252 20269 17255
rect 19260 17224 20269 17252
rect 16669 17187 16727 17193
rect 16669 17153 16681 17187
rect 16715 17153 16727 17187
rect 17034 17184 17040 17196
rect 16995 17156 17040 17184
rect 16669 17147 16727 17153
rect 17034 17144 17040 17156
rect 17092 17144 17098 17196
rect 19061 17187 19119 17193
rect 19061 17153 19073 17187
rect 19107 17153 19119 17187
rect 19061 17147 19119 17153
rect 19076 17116 19104 17147
rect 19150 17144 19156 17196
rect 19208 17184 19214 17196
rect 19260 17193 19288 17224
rect 20257 17221 20269 17224
rect 20303 17221 20315 17255
rect 20257 17215 20315 17221
rect 20349 17255 20407 17261
rect 20349 17221 20361 17255
rect 20395 17252 20407 17255
rect 22066 17252 22094 17292
rect 25961 17289 25973 17292
rect 26007 17289 26019 17323
rect 25961 17283 26019 17289
rect 20395 17224 22094 17252
rect 20395 17221 20407 17224
rect 20349 17215 20407 17221
rect 22738 17212 22744 17264
rect 22796 17252 22802 17264
rect 22796 17224 24992 17252
rect 22796 17212 22802 17224
rect 19245 17187 19303 17193
rect 19245 17184 19257 17187
rect 19208 17156 19257 17184
rect 19208 17144 19214 17156
rect 19245 17153 19257 17156
rect 19291 17153 19303 17187
rect 19245 17147 19303 17153
rect 19337 17187 19395 17193
rect 19337 17153 19349 17187
rect 19383 17153 19395 17187
rect 19337 17147 19395 17153
rect 19429 17187 19487 17193
rect 19429 17153 19441 17187
rect 19475 17153 19487 17187
rect 19429 17147 19487 17153
rect 20073 17187 20131 17193
rect 20073 17153 20085 17187
rect 20119 17184 20131 17187
rect 20162 17184 20168 17196
rect 20119 17156 20168 17184
rect 20119 17153 20131 17156
rect 20073 17147 20131 17153
rect 15212 17088 19104 17116
rect 17034 17008 17040 17060
rect 17092 17048 17098 17060
rect 18049 17051 18107 17057
rect 18049 17048 18061 17051
rect 17092 17020 18061 17048
rect 17092 17008 17098 17020
rect 18049 17017 18061 17020
rect 18095 17017 18107 17051
rect 19352 17048 19380 17147
rect 19444 17116 19472 17147
rect 20162 17144 20168 17156
rect 20220 17144 20226 17196
rect 20441 17187 20499 17193
rect 20441 17153 20453 17187
rect 20487 17153 20499 17187
rect 20441 17147 20499 17153
rect 19518 17116 19524 17128
rect 19444 17088 19524 17116
rect 19518 17076 19524 17088
rect 19576 17116 19582 17128
rect 20456 17116 20484 17147
rect 20898 17144 20904 17196
rect 20956 17184 20962 17196
rect 21085 17187 21143 17193
rect 21085 17184 21097 17187
rect 20956 17156 21097 17184
rect 20956 17144 20962 17156
rect 21085 17153 21097 17156
rect 21131 17153 21143 17187
rect 21085 17147 21143 17153
rect 22094 17144 22100 17196
rect 22152 17184 22158 17196
rect 23492 17193 23520 17224
rect 23477 17187 23535 17193
rect 22152 17156 22197 17184
rect 22152 17144 22158 17156
rect 23477 17153 23489 17187
rect 23523 17153 23535 17187
rect 23750 17184 23756 17196
rect 23711 17156 23756 17184
rect 23477 17147 23535 17153
rect 23750 17144 23756 17156
rect 23808 17144 23814 17196
rect 24964 17193 24992 17224
rect 24949 17187 25007 17193
rect 24949 17153 24961 17187
rect 24995 17153 25007 17187
rect 25222 17184 25228 17196
rect 25183 17156 25228 17184
rect 24949 17147 25007 17153
rect 25222 17144 25228 17156
rect 25280 17144 25286 17196
rect 19576 17088 20484 17116
rect 19576 17076 19582 17088
rect 21450 17076 21456 17128
rect 21508 17116 21514 17128
rect 21821 17119 21879 17125
rect 21821 17116 21833 17119
rect 21508 17088 21833 17116
rect 21508 17076 21514 17088
rect 21821 17085 21833 17088
rect 21867 17085 21879 17119
rect 21821 17079 21879 17085
rect 19352 17020 20760 17048
rect 18049 17011 18107 17017
rect 12618 16940 12624 16992
rect 12676 16980 12682 16992
rect 12805 16983 12863 16989
rect 12805 16980 12817 16983
rect 12676 16952 12817 16980
rect 12676 16940 12682 16952
rect 12805 16949 12817 16952
rect 12851 16949 12863 16983
rect 17218 16980 17224 16992
rect 17179 16952 17224 16980
rect 12805 16943 12863 16949
rect 17218 16940 17224 16952
rect 17276 16940 17282 16992
rect 17865 16983 17923 16989
rect 17865 16949 17877 16983
rect 17911 16980 17923 16983
rect 18138 16980 18144 16992
rect 17911 16952 18144 16980
rect 17911 16949 17923 16952
rect 17865 16943 17923 16949
rect 18138 16940 18144 16952
rect 18196 16940 18202 16992
rect 19426 16940 19432 16992
rect 19484 16980 19490 16992
rect 19613 16983 19671 16989
rect 19613 16980 19625 16983
rect 19484 16952 19625 16980
rect 19484 16940 19490 16952
rect 19613 16949 19625 16952
rect 19659 16949 19671 16983
rect 19613 16943 19671 16949
rect 20254 16940 20260 16992
rect 20312 16980 20318 16992
rect 20625 16983 20683 16989
rect 20625 16980 20637 16983
rect 20312 16952 20637 16980
rect 20312 16940 20318 16952
rect 20625 16949 20637 16952
rect 20671 16949 20683 16983
rect 20732 16980 20760 17020
rect 22756 17020 23060 17048
rect 22756 16980 22784 17020
rect 20732 16952 22784 16980
rect 20625 16943 20683 16949
rect 22830 16940 22836 16992
rect 22888 16980 22894 16992
rect 23032 16980 23060 17020
rect 24489 16983 24547 16989
rect 24489 16980 24501 16983
rect 22888 16952 22933 16980
rect 23032 16952 24501 16980
rect 22888 16940 22894 16952
rect 24489 16949 24501 16952
rect 24535 16949 24547 16983
rect 24489 16943 24547 16949
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 10594 16736 10600 16788
rect 10652 16776 10658 16788
rect 12345 16779 12403 16785
rect 12345 16776 12357 16779
rect 10652 16748 12357 16776
rect 10652 16736 10658 16748
rect 12345 16745 12357 16748
rect 12391 16745 12403 16779
rect 12802 16776 12808 16788
rect 12763 16748 12808 16776
rect 12345 16739 12403 16745
rect 12802 16736 12808 16748
rect 12860 16736 12866 16788
rect 14182 16736 14188 16788
rect 14240 16776 14246 16788
rect 20070 16776 20076 16788
rect 14240 16748 20076 16776
rect 14240 16736 14246 16748
rect 12710 16708 12716 16720
rect 12544 16680 12716 16708
rect 9398 16600 9404 16652
rect 9456 16640 9462 16652
rect 9861 16643 9919 16649
rect 9861 16640 9873 16643
rect 9456 16612 9873 16640
rect 9456 16600 9462 16612
rect 9861 16609 9873 16612
rect 9907 16609 9919 16643
rect 9861 16603 9919 16609
rect 12544 16581 12572 16680
rect 12710 16668 12716 16680
rect 12768 16708 12774 16720
rect 14093 16711 14151 16717
rect 14093 16708 14105 16711
rect 12768 16680 14105 16708
rect 12768 16668 12774 16680
rect 14093 16677 14105 16680
rect 14139 16677 14151 16711
rect 14734 16708 14740 16720
rect 14695 16680 14740 16708
rect 14093 16671 14151 16677
rect 14734 16668 14740 16680
rect 14792 16668 14798 16720
rect 13078 16600 13084 16652
rect 13136 16640 13142 16652
rect 15488 16649 15516 16748
rect 20070 16736 20076 16748
rect 20128 16776 20134 16788
rect 20128 16748 25176 16776
rect 20128 16736 20134 16748
rect 16853 16711 16911 16717
rect 16853 16677 16865 16711
rect 16899 16708 16911 16711
rect 16942 16708 16948 16720
rect 16899 16680 16948 16708
rect 16899 16677 16911 16680
rect 16853 16671 16911 16677
rect 16942 16668 16948 16680
rect 17000 16668 17006 16720
rect 18049 16711 18107 16717
rect 18049 16677 18061 16711
rect 18095 16708 18107 16711
rect 18230 16708 18236 16720
rect 18095 16680 18236 16708
rect 18095 16677 18107 16680
rect 18049 16671 18107 16677
rect 18230 16668 18236 16680
rect 18288 16668 18294 16720
rect 20349 16711 20407 16717
rect 20349 16677 20361 16711
rect 20395 16708 20407 16711
rect 20990 16708 20996 16720
rect 20395 16680 20996 16708
rect 20395 16677 20407 16680
rect 20349 16671 20407 16677
rect 20990 16668 20996 16680
rect 21048 16668 21054 16720
rect 25148 16649 25176 16748
rect 15473 16643 15531 16649
rect 13136 16612 14320 16640
rect 13136 16600 13142 16612
rect 12529 16575 12587 16581
rect 12529 16541 12541 16575
rect 12575 16541 12587 16575
rect 12529 16535 12587 16541
rect 12618 16532 12624 16584
rect 12676 16572 12682 16584
rect 12894 16572 12900 16584
rect 12676 16544 12721 16572
rect 12855 16544 12900 16572
rect 12676 16532 12682 16544
rect 12894 16532 12900 16544
rect 12952 16532 12958 16584
rect 13538 16572 13544 16584
rect 13499 16544 13544 16572
rect 13538 16532 13544 16544
rect 13596 16532 13602 16584
rect 14090 16572 14096 16584
rect 14051 16544 14096 16572
rect 14090 16532 14096 16544
rect 14148 16532 14154 16584
rect 14292 16581 14320 16612
rect 15473 16609 15485 16643
rect 15519 16609 15531 16643
rect 15473 16603 15531 16609
rect 25133 16643 25191 16649
rect 25133 16609 25145 16643
rect 25179 16609 25191 16643
rect 25133 16603 25191 16609
rect 14277 16575 14335 16581
rect 14277 16541 14289 16575
rect 14323 16541 14335 16575
rect 14918 16572 14924 16584
rect 14879 16544 14924 16572
rect 14277 16535 14335 16541
rect 14918 16532 14924 16544
rect 14976 16532 14982 16584
rect 15740 16575 15798 16581
rect 15740 16541 15752 16575
rect 15786 16572 15798 16575
rect 17218 16572 17224 16584
rect 15786 16544 17224 16572
rect 15786 16541 15798 16544
rect 15740 16535 15798 16541
rect 17218 16532 17224 16544
rect 17276 16532 17282 16584
rect 17862 16572 17868 16584
rect 17823 16544 17868 16572
rect 17862 16532 17868 16544
rect 17920 16532 17926 16584
rect 18690 16572 18696 16584
rect 18651 16544 18696 16572
rect 18690 16532 18696 16544
rect 18748 16532 18754 16584
rect 19334 16572 19340 16584
rect 19295 16544 19340 16572
rect 19334 16532 19340 16544
rect 19392 16532 19398 16584
rect 19613 16575 19671 16581
rect 19613 16541 19625 16575
rect 19659 16541 19671 16575
rect 21450 16572 21456 16584
rect 21411 16544 21456 16572
rect 19613 16535 19671 16541
rect 9582 16464 9588 16516
rect 9640 16504 9646 16516
rect 10106 16507 10164 16513
rect 10106 16504 10118 16507
rect 9640 16476 10118 16504
rect 9640 16464 9646 16476
rect 10106 16473 10118 16476
rect 10152 16473 10164 16507
rect 10106 16467 10164 16473
rect 19150 16464 19156 16516
rect 19208 16504 19214 16516
rect 19628 16504 19656 16535
rect 21450 16532 21456 16544
rect 21508 16532 21514 16584
rect 21729 16575 21787 16581
rect 21729 16541 21741 16575
rect 21775 16572 21787 16575
rect 23014 16572 23020 16584
rect 21775 16544 23020 16572
rect 21775 16541 21787 16544
rect 21729 16535 21787 16541
rect 23014 16532 23020 16544
rect 23072 16532 23078 16584
rect 23385 16575 23443 16581
rect 23385 16541 23397 16575
rect 23431 16572 23443 16575
rect 23750 16572 23756 16584
rect 23431 16544 23756 16572
rect 23431 16541 23443 16544
rect 23385 16535 23443 16541
rect 23750 16532 23756 16544
rect 23808 16532 23814 16584
rect 25406 16572 25412 16584
rect 25367 16544 25412 16572
rect 25406 16532 25412 16544
rect 25464 16532 25470 16584
rect 19208 16476 19656 16504
rect 19208 16464 19214 16476
rect 11241 16439 11299 16445
rect 11241 16405 11253 16439
rect 11287 16436 11299 16439
rect 11790 16436 11796 16448
rect 11287 16408 11796 16436
rect 11287 16405 11299 16408
rect 11241 16399 11299 16405
rect 11790 16396 11796 16408
rect 11848 16396 11854 16448
rect 13354 16436 13360 16448
rect 13315 16408 13360 16436
rect 13354 16396 13360 16408
rect 13412 16396 13418 16448
rect 18509 16439 18567 16445
rect 18509 16405 18521 16439
rect 18555 16436 18567 16439
rect 18690 16436 18696 16448
rect 18555 16408 18696 16436
rect 18555 16405 18567 16408
rect 18509 16399 18567 16405
rect 18690 16396 18696 16408
rect 18748 16396 18754 16448
rect 22462 16436 22468 16448
rect 22423 16408 22468 16436
rect 22462 16396 22468 16408
rect 22520 16396 22526 16448
rect 23198 16436 23204 16448
rect 23159 16408 23204 16436
rect 23198 16396 23204 16408
rect 23256 16396 23262 16448
rect 23474 16396 23480 16448
rect 23532 16436 23538 16448
rect 24394 16436 24400 16448
rect 23532 16408 24400 16436
rect 23532 16396 23538 16408
rect 24394 16396 24400 16408
rect 24452 16396 24458 16448
rect 25682 16396 25688 16448
rect 25740 16436 25746 16448
rect 26513 16439 26571 16445
rect 26513 16436 26525 16439
rect 25740 16408 26525 16436
rect 25740 16396 25746 16408
rect 26513 16405 26525 16408
rect 26559 16405 26571 16439
rect 26513 16399 26571 16405
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 11977 16235 12035 16241
rect 11977 16201 11989 16235
rect 12023 16232 12035 16235
rect 12618 16232 12624 16244
rect 12023 16204 12624 16232
rect 12023 16201 12035 16204
rect 11977 16195 12035 16201
rect 12618 16192 12624 16204
rect 12676 16192 12682 16244
rect 13817 16235 13875 16241
rect 13817 16201 13829 16235
rect 13863 16232 13875 16235
rect 14090 16232 14096 16244
rect 13863 16204 14096 16232
rect 13863 16201 13875 16204
rect 13817 16195 13875 16201
rect 14090 16192 14096 16204
rect 14148 16192 14154 16244
rect 16482 16232 16488 16244
rect 16443 16204 16488 16232
rect 16482 16192 16488 16204
rect 16540 16192 16546 16244
rect 18509 16235 18567 16241
rect 18509 16201 18521 16235
rect 18555 16232 18567 16235
rect 19334 16232 19340 16244
rect 18555 16204 19340 16232
rect 18555 16201 18567 16204
rect 18509 16195 18567 16201
rect 19334 16192 19340 16204
rect 19392 16192 19398 16244
rect 22554 16192 22560 16244
rect 22612 16232 22618 16244
rect 22833 16235 22891 16241
rect 22833 16232 22845 16235
rect 22612 16204 22845 16232
rect 22612 16192 22618 16204
rect 22833 16201 22845 16204
rect 22879 16201 22891 16235
rect 24949 16235 25007 16241
rect 24949 16232 24961 16235
rect 22833 16195 22891 16201
rect 23124 16204 24961 16232
rect 9398 16164 9404 16176
rect 8588 16136 9404 16164
rect 8588 16108 8616 16136
rect 9398 16124 9404 16136
rect 9456 16124 9462 16176
rect 12704 16167 12762 16173
rect 12704 16133 12716 16167
rect 12750 16164 12762 16167
rect 13354 16164 13360 16176
rect 12750 16136 13360 16164
rect 12750 16133 12762 16136
rect 12704 16127 12762 16133
rect 13354 16124 13360 16136
rect 13412 16124 13418 16176
rect 22741 16167 22799 16173
rect 17788 16136 22094 16164
rect 7929 16099 7987 16105
rect 7929 16065 7941 16099
rect 7975 16096 7987 16099
rect 8294 16096 8300 16108
rect 7975 16068 8300 16096
rect 7975 16065 7987 16068
rect 7929 16059 7987 16065
rect 8294 16056 8300 16068
rect 8352 16056 8358 16108
rect 8570 16096 8576 16108
rect 8483 16068 8576 16096
rect 8570 16056 8576 16068
rect 8628 16056 8634 16108
rect 8846 16105 8852 16108
rect 8840 16059 8852 16105
rect 8904 16096 8910 16108
rect 12437 16099 12495 16105
rect 8904 16068 8940 16096
rect 8846 16056 8852 16059
rect 8904 16056 8910 16068
rect 12437 16065 12449 16099
rect 12483 16096 12495 16099
rect 13170 16096 13176 16108
rect 12483 16068 13176 16096
rect 12483 16065 12495 16068
rect 12437 16059 12495 16065
rect 13170 16056 13176 16068
rect 13228 16056 13234 16108
rect 14182 16056 14188 16108
rect 14240 16096 14246 16108
rect 17788 16105 17816 16136
rect 14461 16099 14519 16105
rect 14461 16096 14473 16099
rect 14240 16068 14473 16096
rect 14240 16056 14246 16068
rect 14461 16065 14473 16068
rect 14507 16065 14519 16099
rect 14461 16059 14519 16065
rect 14728 16099 14786 16105
rect 14728 16065 14740 16099
rect 14774 16096 14786 16099
rect 17313 16099 17371 16105
rect 14774 16068 16160 16096
rect 14774 16065 14786 16068
rect 14728 16059 14786 16065
rect 11517 16031 11575 16037
rect 11517 15997 11529 16031
rect 11563 16028 11575 16031
rect 12250 16028 12256 16040
rect 11563 16000 12256 16028
rect 11563 15997 11575 16000
rect 11517 15991 11575 15997
rect 12250 15988 12256 16000
rect 12308 15988 12314 16040
rect 16025 16031 16083 16037
rect 16025 15997 16037 16031
rect 16071 15997 16083 16031
rect 16025 15991 16083 15997
rect 11790 15960 11796 15972
rect 11751 15932 11796 15960
rect 11790 15920 11796 15932
rect 11848 15920 11854 15972
rect 15841 15963 15899 15969
rect 15841 15929 15853 15963
rect 15887 15960 15899 15963
rect 16040 15960 16068 15991
rect 15887 15932 16068 15960
rect 16132 15960 16160 16068
rect 17313 16065 17325 16099
rect 17359 16096 17371 16099
rect 17773 16099 17831 16105
rect 17773 16096 17785 16099
rect 17359 16068 17785 16096
rect 17359 16065 17371 16068
rect 17313 16059 17371 16065
rect 17773 16065 17785 16068
rect 17819 16065 17831 16099
rect 18690 16096 18696 16108
rect 18651 16068 18696 16096
rect 17773 16059 17831 16065
rect 18690 16056 18696 16068
rect 18748 16056 18754 16108
rect 19334 16056 19340 16108
rect 19392 16096 19398 16108
rect 19429 16099 19487 16105
rect 19429 16096 19441 16099
rect 19392 16068 19441 16096
rect 19392 16056 19398 16068
rect 19429 16065 19441 16068
rect 19475 16065 19487 16099
rect 20254 16096 20260 16108
rect 20215 16068 20260 16096
rect 19429 16059 19487 16065
rect 20254 16056 20260 16068
rect 20312 16056 20318 16108
rect 22066 16096 22094 16136
rect 22741 16133 22753 16167
rect 22787 16164 22799 16167
rect 23124 16164 23152 16204
rect 24949 16201 24961 16204
rect 24995 16232 25007 16235
rect 25038 16232 25044 16244
rect 24995 16204 25044 16232
rect 24995 16201 25007 16204
rect 24949 16195 25007 16201
rect 25038 16192 25044 16204
rect 25096 16192 25102 16244
rect 25406 16192 25412 16244
rect 25464 16232 25470 16244
rect 25501 16235 25559 16241
rect 25501 16232 25513 16235
rect 25464 16204 25513 16232
rect 25464 16192 25470 16204
rect 25501 16201 25513 16204
rect 25547 16201 25559 16235
rect 25501 16195 25559 16201
rect 22787 16136 23152 16164
rect 22787 16133 22799 16136
rect 22741 16127 22799 16133
rect 23198 16124 23204 16176
rect 23256 16164 23262 16176
rect 23814 16167 23872 16173
rect 23814 16164 23826 16167
rect 23256 16136 23826 16164
rect 23256 16124 23262 16136
rect 23814 16133 23826 16136
rect 23860 16133 23872 16167
rect 23814 16127 23872 16133
rect 24412 16136 25636 16164
rect 23474 16096 23480 16108
rect 22066 16068 23480 16096
rect 23474 16056 23480 16068
rect 23532 16056 23538 16108
rect 23569 16099 23627 16105
rect 23569 16065 23581 16099
rect 23615 16096 23627 16099
rect 24412 16096 24440 16136
rect 23615 16068 24440 16096
rect 25409 16099 25467 16105
rect 23615 16065 23627 16068
rect 23569 16059 23627 16065
rect 25409 16065 25421 16099
rect 25455 16096 25467 16099
rect 25498 16096 25504 16108
rect 25455 16068 25504 16096
rect 25455 16065 25467 16068
rect 25409 16059 25467 16065
rect 25498 16056 25504 16068
rect 25556 16056 25562 16108
rect 25608 16105 25636 16136
rect 25593 16099 25651 16105
rect 25593 16065 25605 16099
rect 25639 16096 25651 16099
rect 25682 16096 25688 16108
rect 25639 16068 25688 16096
rect 25639 16065 25651 16068
rect 25593 16059 25651 16065
rect 25682 16056 25688 16068
rect 25740 16056 25746 16108
rect 26050 16096 26056 16108
rect 26011 16068 26056 16096
rect 26050 16056 26056 16068
rect 26108 16056 26114 16108
rect 26237 16099 26295 16105
rect 26237 16065 26249 16099
rect 26283 16065 26295 16099
rect 26237 16059 26295 16065
rect 17957 16031 18015 16037
rect 17957 15997 17969 16031
rect 18003 16028 18015 16031
rect 18046 16028 18052 16040
rect 18003 16000 18052 16028
rect 18003 15997 18015 16000
rect 17957 15991 18015 15997
rect 18046 15988 18052 16000
rect 18104 15988 18110 16040
rect 19150 15988 19156 16040
rect 19208 16028 19214 16040
rect 19981 16031 20039 16037
rect 19981 16028 19993 16031
rect 19208 16000 19993 16028
rect 19208 15988 19214 16000
rect 19981 15997 19993 16000
rect 20027 15997 20039 16031
rect 22922 16028 22928 16040
rect 22883 16000 22928 16028
rect 19981 15991 20039 15997
rect 22922 15988 22928 16000
rect 22980 15988 22986 16040
rect 25516 16028 25544 16056
rect 26252 16028 26280 16059
rect 25516 16000 26280 16028
rect 16301 15963 16359 15969
rect 16301 15960 16313 15963
rect 16132 15932 16313 15960
rect 15887 15929 15899 15932
rect 15841 15923 15899 15929
rect 16301 15929 16313 15932
rect 16347 15960 16359 15963
rect 16390 15960 16396 15972
rect 16347 15932 16396 15960
rect 16347 15929 16359 15932
rect 16301 15923 16359 15929
rect 16390 15920 16396 15932
rect 16448 15920 16454 15972
rect 18874 15920 18880 15972
rect 18932 15960 18938 15972
rect 19245 15963 19303 15969
rect 19245 15960 19257 15963
rect 18932 15932 19257 15960
rect 18932 15920 18938 15932
rect 19245 15929 19257 15932
rect 19291 15929 19303 15963
rect 19245 15923 19303 15929
rect 7742 15892 7748 15904
rect 7703 15864 7748 15892
rect 7742 15852 7748 15864
rect 7800 15852 7806 15904
rect 9950 15892 9956 15904
rect 9911 15864 9956 15892
rect 9950 15852 9956 15864
rect 10008 15852 10014 15904
rect 17586 15892 17592 15904
rect 17547 15864 17592 15892
rect 17586 15852 17592 15864
rect 17644 15852 17650 15904
rect 20993 15895 21051 15901
rect 20993 15861 21005 15895
rect 21039 15892 21051 15895
rect 22094 15892 22100 15904
rect 21039 15864 22100 15892
rect 21039 15861 21051 15864
rect 20993 15855 21051 15861
rect 22094 15852 22100 15864
rect 22152 15852 22158 15904
rect 22373 15895 22431 15901
rect 22373 15861 22385 15895
rect 22419 15892 22431 15895
rect 23566 15892 23572 15904
rect 22419 15864 23572 15892
rect 22419 15861 22431 15864
rect 22373 15855 22431 15861
rect 23566 15852 23572 15864
rect 23624 15852 23630 15904
rect 26053 15895 26111 15901
rect 26053 15861 26065 15895
rect 26099 15892 26111 15895
rect 26234 15892 26240 15904
rect 26099 15864 26240 15892
rect 26099 15861 26111 15864
rect 26053 15855 26111 15861
rect 26234 15852 26240 15864
rect 26292 15852 26298 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 8570 15688 8576 15700
rect 7024 15660 8576 15688
rect 7024 15564 7052 15660
rect 8570 15648 8576 15660
rect 8628 15648 8634 15700
rect 8846 15648 8852 15700
rect 8904 15688 8910 15700
rect 8941 15691 8999 15697
rect 8941 15688 8953 15691
rect 8904 15660 8953 15688
rect 8904 15648 8910 15660
rect 8941 15657 8953 15660
rect 8987 15657 8999 15691
rect 9582 15688 9588 15700
rect 9543 15660 9588 15688
rect 8941 15651 8999 15657
rect 9582 15648 9588 15660
rect 9640 15648 9646 15700
rect 12529 15691 12587 15697
rect 12529 15657 12541 15691
rect 12575 15688 12587 15691
rect 12894 15688 12900 15700
rect 12575 15660 12900 15688
rect 12575 15657 12587 15660
rect 12529 15651 12587 15657
rect 12894 15648 12900 15660
rect 12952 15648 12958 15700
rect 13357 15691 13415 15697
rect 13357 15657 13369 15691
rect 13403 15688 13415 15691
rect 13538 15688 13544 15700
rect 13403 15660 13544 15688
rect 13403 15657 13415 15660
rect 13357 15651 13415 15657
rect 13538 15648 13544 15660
rect 13596 15648 13602 15700
rect 18230 15688 18236 15700
rect 17788 15660 18236 15688
rect 12250 15580 12256 15632
rect 12308 15620 12314 15632
rect 12345 15623 12403 15629
rect 12345 15620 12357 15623
rect 12308 15592 12357 15620
rect 12308 15580 12314 15592
rect 12345 15589 12357 15592
rect 12391 15589 12403 15623
rect 17788 15620 17816 15660
rect 18230 15648 18236 15660
rect 18288 15648 18294 15700
rect 21450 15688 21456 15700
rect 19260 15660 21456 15688
rect 12345 15583 12403 15589
rect 17696 15592 17816 15620
rect 18248 15620 18276 15648
rect 19150 15620 19156 15632
rect 18248 15592 19156 15620
rect 7006 15552 7012 15564
rect 6919 15524 7012 15552
rect 7006 15512 7012 15524
rect 7064 15512 7070 15564
rect 9950 15552 9956 15564
rect 9911 15524 9956 15552
rect 9950 15512 9956 15524
rect 10008 15512 10014 15564
rect 10045 15555 10103 15561
rect 10045 15521 10057 15555
rect 10091 15552 10103 15555
rect 10597 15555 10655 15561
rect 10597 15552 10609 15555
rect 10091 15524 10609 15552
rect 10091 15521 10103 15524
rect 10045 15515 10103 15521
rect 10597 15521 10609 15524
rect 10643 15521 10655 15555
rect 11790 15552 11796 15564
rect 10597 15515 10655 15521
rect 11072 15524 11796 15552
rect 7276 15487 7334 15493
rect 7276 15453 7288 15487
rect 7322 15484 7334 15487
rect 7742 15484 7748 15496
rect 7322 15456 7748 15484
rect 7322 15453 7334 15456
rect 7276 15447 7334 15453
rect 7742 15444 7748 15456
rect 7800 15444 7806 15496
rect 9122 15484 9128 15496
rect 9083 15456 9128 15484
rect 9122 15444 9128 15456
rect 9180 15444 9186 15496
rect 9766 15484 9772 15496
rect 9727 15456 9772 15484
rect 9766 15444 9772 15456
rect 9824 15444 9830 15496
rect 9858 15444 9864 15496
rect 9916 15484 9922 15496
rect 10870 15484 10876 15496
rect 9916 15456 9961 15484
rect 10831 15456 10876 15484
rect 9916 15444 9922 15456
rect 10870 15444 10876 15456
rect 10928 15444 10934 15496
rect 11072 15493 11100 15524
rect 11790 15512 11796 15524
rect 11848 15552 11854 15564
rect 17696 15561 17724 15592
rect 19150 15580 19156 15592
rect 19208 15620 19214 15632
rect 19260 15620 19288 15660
rect 19208 15592 19288 15620
rect 19208 15580 19214 15592
rect 19260 15561 19288 15592
rect 20732 15561 20760 15660
rect 21450 15648 21456 15660
rect 21508 15648 21514 15700
rect 23750 15688 23756 15700
rect 23711 15660 23756 15688
rect 23750 15648 23756 15660
rect 23808 15648 23814 15700
rect 25038 15688 25044 15700
rect 24999 15660 25044 15688
rect 25038 15648 25044 15660
rect 25096 15648 25102 15700
rect 25961 15691 26019 15697
rect 25961 15657 25973 15691
rect 26007 15688 26019 15691
rect 26050 15688 26056 15700
rect 26007 15660 26056 15688
rect 26007 15657 26019 15660
rect 25961 15651 26019 15657
rect 25976 15620 26004 15651
rect 26050 15648 26056 15660
rect 26108 15648 26114 15700
rect 25332 15592 26004 15620
rect 12069 15555 12127 15561
rect 12069 15552 12081 15555
rect 11848 15524 12081 15552
rect 11848 15512 11854 15524
rect 12069 15521 12081 15524
rect 12115 15552 12127 15555
rect 12989 15555 13047 15561
rect 12989 15552 13001 15555
rect 12115 15524 13001 15552
rect 12115 15521 12127 15524
rect 12069 15515 12127 15521
rect 12989 15521 13001 15524
rect 13035 15521 13047 15555
rect 12989 15515 13047 15521
rect 17681 15555 17739 15561
rect 17681 15521 17693 15555
rect 17727 15521 17739 15555
rect 17681 15515 17739 15521
rect 19245 15555 19303 15561
rect 19245 15521 19257 15555
rect 19291 15521 19303 15555
rect 19245 15515 19303 15521
rect 20717 15555 20775 15561
rect 20717 15521 20729 15555
rect 20763 15521 20775 15555
rect 20717 15515 20775 15521
rect 22462 15512 22468 15564
rect 22520 15552 22526 15564
rect 22649 15555 22707 15561
rect 22649 15552 22661 15555
rect 22520 15524 22661 15552
rect 22520 15512 22526 15524
rect 22649 15521 22661 15524
rect 22695 15521 22707 15555
rect 22649 15515 22707 15521
rect 22833 15555 22891 15561
rect 22833 15521 22845 15555
rect 22879 15552 22891 15555
rect 22922 15552 22928 15564
rect 22879 15524 22928 15552
rect 22879 15521 22891 15524
rect 22833 15515 22891 15521
rect 10965 15487 11023 15493
rect 10965 15453 10977 15487
rect 11011 15453 11023 15487
rect 10965 15447 11023 15453
rect 11057 15487 11115 15493
rect 11057 15453 11069 15487
rect 11103 15453 11115 15487
rect 11057 15447 11115 15453
rect 11241 15487 11299 15493
rect 11241 15453 11253 15487
rect 11287 15484 11299 15487
rect 11330 15484 11336 15496
rect 11287 15456 11336 15484
rect 11287 15453 11299 15456
rect 11241 15447 11299 15453
rect 10134 15376 10140 15428
rect 10192 15416 10198 15428
rect 10980 15416 11008 15447
rect 11330 15444 11336 15456
rect 11388 15444 11394 15496
rect 13173 15487 13231 15493
rect 13173 15453 13185 15487
rect 13219 15484 13231 15487
rect 13446 15484 13452 15496
rect 13219 15456 13452 15484
rect 13219 15453 13231 15456
rect 13173 15447 13231 15453
rect 13446 15444 13452 15456
rect 13504 15444 13510 15496
rect 15010 15444 15016 15496
rect 15068 15484 15074 15496
rect 15565 15487 15623 15493
rect 15565 15484 15577 15487
rect 15068 15456 15577 15484
rect 15068 15444 15074 15456
rect 15565 15453 15577 15456
rect 15611 15453 15623 15487
rect 17954 15484 17960 15496
rect 17915 15456 17960 15484
rect 15565 15447 15623 15453
rect 17954 15444 17960 15456
rect 18012 15444 18018 15496
rect 19426 15444 19432 15496
rect 19484 15484 19490 15496
rect 19521 15487 19579 15493
rect 19521 15484 19533 15487
rect 19484 15456 19533 15484
rect 19484 15444 19490 15456
rect 19521 15453 19533 15456
rect 19567 15453 19579 15487
rect 19521 15447 19579 15453
rect 20993 15487 21051 15493
rect 20993 15453 21005 15487
rect 21039 15484 21051 15487
rect 21082 15484 21088 15496
rect 21039 15456 21088 15484
rect 21039 15453 21051 15456
rect 20993 15447 21051 15453
rect 21082 15444 21088 15456
rect 21140 15444 21146 15496
rect 22370 15444 22376 15496
rect 22428 15484 22434 15496
rect 22848 15484 22876 15515
rect 22922 15512 22928 15524
rect 22980 15512 22986 15564
rect 22428 15456 22876 15484
rect 23385 15487 23443 15493
rect 22428 15444 22434 15456
rect 23385 15453 23397 15487
rect 23431 15453 23443 15487
rect 23566 15484 23572 15496
rect 23527 15456 23572 15484
rect 23385 15447 23443 15453
rect 10192 15388 11008 15416
rect 15832 15419 15890 15425
rect 10192 15376 10198 15388
rect 15832 15385 15844 15419
rect 15878 15416 15890 15419
rect 16666 15416 16672 15428
rect 15878 15388 16672 15416
rect 15878 15385 15890 15388
rect 15832 15379 15890 15385
rect 16666 15376 16672 15388
rect 16724 15376 16730 15428
rect 22738 15376 22744 15428
rect 22796 15416 22802 15428
rect 23400 15416 23428 15447
rect 23566 15444 23572 15456
rect 23624 15444 23630 15496
rect 24949 15487 25007 15493
rect 24949 15453 24961 15487
rect 24995 15484 25007 15487
rect 25332 15484 25360 15592
rect 26145 15555 26203 15561
rect 26145 15552 26157 15555
rect 24995 15456 25360 15484
rect 25424 15524 26157 15552
rect 24995 15453 25007 15456
rect 24949 15447 25007 15453
rect 22796 15388 23428 15416
rect 22796 15376 22802 15388
rect 8386 15348 8392 15360
rect 8299 15320 8392 15348
rect 8386 15308 8392 15320
rect 8444 15348 8450 15360
rect 9582 15348 9588 15360
rect 8444 15320 9588 15348
rect 8444 15308 8450 15320
rect 9582 15308 9588 15320
rect 9640 15308 9646 15360
rect 15194 15308 15200 15360
rect 15252 15348 15258 15360
rect 16945 15351 17003 15357
rect 16945 15348 16957 15351
rect 15252 15320 16957 15348
rect 15252 15308 15258 15320
rect 16945 15317 16957 15320
rect 16991 15317 17003 15351
rect 16945 15311 17003 15317
rect 18414 15308 18420 15360
rect 18472 15348 18478 15360
rect 18693 15351 18751 15357
rect 18693 15348 18705 15351
rect 18472 15320 18705 15348
rect 18472 15308 18478 15320
rect 18693 15317 18705 15320
rect 18739 15317 18751 15351
rect 20254 15348 20260 15360
rect 20215 15320 20260 15348
rect 18693 15311 18751 15317
rect 20254 15308 20260 15320
rect 20312 15308 20318 15360
rect 20806 15308 20812 15360
rect 20864 15348 20870 15360
rect 21729 15351 21787 15357
rect 21729 15348 21741 15351
rect 20864 15320 21741 15348
rect 20864 15308 20870 15320
rect 21729 15317 21741 15320
rect 21775 15317 21787 15351
rect 21729 15311 21787 15317
rect 22189 15351 22247 15357
rect 22189 15317 22201 15351
rect 22235 15348 22247 15351
rect 22462 15348 22468 15360
rect 22235 15320 22468 15348
rect 22235 15317 22247 15320
rect 22189 15311 22247 15317
rect 22462 15308 22468 15320
rect 22520 15308 22526 15360
rect 22557 15351 22615 15357
rect 22557 15317 22569 15351
rect 22603 15348 22615 15351
rect 23934 15348 23940 15360
rect 22603 15320 23940 15348
rect 22603 15317 22615 15320
rect 22557 15311 22615 15317
rect 23934 15308 23940 15320
rect 23992 15308 23998 15360
rect 25314 15308 25320 15360
rect 25372 15348 25378 15360
rect 25424 15357 25452 15524
rect 26145 15521 26157 15524
rect 26191 15521 26203 15555
rect 26145 15515 26203 15521
rect 25498 15444 25504 15496
rect 25556 15484 25562 15496
rect 25869 15487 25927 15493
rect 25869 15484 25881 15487
rect 25556 15456 25881 15484
rect 25556 15444 25562 15456
rect 25869 15453 25881 15456
rect 25915 15453 25927 15487
rect 25869 15447 25927 15453
rect 25409 15351 25467 15357
rect 25409 15348 25421 15351
rect 25372 15320 25421 15348
rect 25372 15308 25378 15320
rect 25409 15317 25421 15320
rect 25455 15317 25467 15351
rect 25409 15311 25467 15317
rect 25498 15308 25504 15360
rect 25556 15348 25562 15360
rect 26145 15351 26203 15357
rect 26145 15348 26157 15351
rect 25556 15320 26157 15348
rect 25556 15308 25562 15320
rect 26145 15317 26157 15320
rect 26191 15317 26203 15351
rect 26145 15311 26203 15317
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 8294 15144 8300 15156
rect 8255 15116 8300 15144
rect 8294 15104 8300 15116
rect 8352 15104 8358 15156
rect 9122 15144 9128 15156
rect 9083 15116 9128 15144
rect 9122 15104 9128 15116
rect 9180 15104 9186 15156
rect 12529 15147 12587 15153
rect 12529 15113 12541 15147
rect 12575 15113 12587 15147
rect 16666 15144 16672 15156
rect 16627 15116 16672 15144
rect 12529 15107 12587 15113
rect 7469 15079 7527 15085
rect 7469 15076 7481 15079
rect 6656 15048 7481 15076
rect 6656 15017 6684 15048
rect 7469 15045 7481 15048
rect 7515 15045 7527 15079
rect 8386 15076 8392 15088
rect 7469 15039 7527 15045
rect 8036 15048 8392 15076
rect 6641 15011 6699 15017
rect 6641 14977 6653 15011
rect 6687 14977 6699 15011
rect 6641 14971 6699 14977
rect 7285 15011 7343 15017
rect 7285 14977 7297 15011
rect 7331 15008 7343 15011
rect 8036 15008 8064 15048
rect 8386 15036 8392 15048
rect 8444 15036 8450 15088
rect 9950 15076 9956 15088
rect 8864 15048 9956 15076
rect 7331 14980 8064 15008
rect 8113 15011 8171 15017
rect 7331 14977 7343 14980
rect 7285 14971 7343 14977
rect 8113 14977 8125 15011
rect 8159 15008 8171 15011
rect 8864 15008 8892 15048
rect 9950 15036 9956 15048
rect 10008 15036 10014 15088
rect 12434 15076 12440 15088
rect 11624 15048 12440 15076
rect 8159 14980 8892 15008
rect 8941 15011 8999 15017
rect 8159 14977 8171 14980
rect 8113 14971 8171 14977
rect 8941 14977 8953 15011
rect 8987 14977 8999 15011
rect 8941 14971 8999 14977
rect 7101 14943 7159 14949
rect 7101 14909 7113 14943
rect 7147 14940 7159 14943
rect 7929 14943 7987 14949
rect 7929 14940 7941 14943
rect 7147 14912 7941 14940
rect 7147 14909 7159 14912
rect 7101 14903 7159 14909
rect 7929 14909 7941 14912
rect 7975 14940 7987 14943
rect 8018 14940 8024 14952
rect 7975 14912 8024 14940
rect 7975 14909 7987 14912
rect 7929 14903 7987 14909
rect 8018 14900 8024 14912
rect 8076 14940 8082 14952
rect 8757 14943 8815 14949
rect 8757 14940 8769 14943
rect 8076 14912 8769 14940
rect 8076 14900 8082 14912
rect 8757 14909 8769 14912
rect 8803 14909 8815 14943
rect 8757 14903 8815 14909
rect 6457 14807 6515 14813
rect 6457 14773 6469 14807
rect 6503 14804 6515 14807
rect 6914 14804 6920 14816
rect 6503 14776 6920 14804
rect 6503 14773 6515 14776
rect 6457 14767 6515 14773
rect 6914 14764 6920 14776
rect 6972 14764 6978 14816
rect 8956 14804 8984 14971
rect 9398 14968 9404 15020
rect 9456 15008 9462 15020
rect 9858 15017 9864 15020
rect 9585 15011 9643 15017
rect 9585 15008 9597 15011
rect 9456 14980 9597 15008
rect 9456 14968 9462 14980
rect 9585 14977 9597 14980
rect 9631 14977 9643 15011
rect 9852 15008 9864 15017
rect 9771 14980 9864 15008
rect 9585 14971 9643 14977
rect 9852 14971 9864 14980
rect 9916 15008 9922 15020
rect 10226 15008 10232 15020
rect 9916 14980 10232 15008
rect 9858 14968 9864 14971
rect 9916 14968 9922 14980
rect 10226 14968 10232 14980
rect 10284 14968 10290 15020
rect 11624 15017 11652 15048
rect 12434 15036 12440 15048
rect 12492 15036 12498 15088
rect 12544 15076 12572 15107
rect 16666 15104 16672 15116
rect 16724 15104 16730 15156
rect 21913 15147 21971 15153
rect 21913 15113 21925 15147
rect 21959 15144 21971 15147
rect 23934 15144 23940 15156
rect 21959 15116 22094 15144
rect 23895 15116 23940 15144
rect 21959 15113 21971 15116
rect 21913 15107 21971 15113
rect 13418 15079 13476 15085
rect 13418 15076 13430 15079
rect 12544 15048 13430 15076
rect 13418 15045 13430 15048
rect 13464 15045 13476 15079
rect 13418 15039 13476 15045
rect 18230 15036 18236 15088
rect 18288 15036 18294 15088
rect 20990 15076 20996 15088
rect 20951 15048 20996 15076
rect 20990 15036 20996 15048
rect 21048 15036 21054 15088
rect 22066 15076 22094 15116
rect 23934 15104 23940 15116
rect 23992 15104 23998 15156
rect 25682 15104 25688 15156
rect 25740 15104 25746 15156
rect 22802 15079 22860 15085
rect 22802 15076 22814 15079
rect 22066 15048 22814 15076
rect 22802 15045 22814 15048
rect 22848 15045 22860 15079
rect 25700 15076 25728 15104
rect 22802 15039 22860 15045
rect 24412 15048 25728 15076
rect 11609 15011 11667 15017
rect 11609 14977 11621 15011
rect 11655 14977 11667 15011
rect 11609 14971 11667 14977
rect 11701 15011 11759 15017
rect 11701 14977 11713 15011
rect 11747 14977 11759 15011
rect 12710 15008 12716 15020
rect 12671 14980 12716 15008
rect 11701 14971 11759 14977
rect 10594 14900 10600 14952
rect 10652 14940 10658 14952
rect 11716 14940 11744 14971
rect 12710 14968 12716 14980
rect 12768 14968 12774 15020
rect 15194 15008 15200 15020
rect 13096 14980 15200 15008
rect 13096 14940 13124 14980
rect 15194 14968 15200 14980
rect 15252 14968 15258 15020
rect 16853 15011 16911 15017
rect 16853 14977 16865 15011
rect 16899 15008 16911 15011
rect 17586 15008 17592 15020
rect 16899 14980 17592 15008
rect 16899 14977 16911 14980
rect 16853 14971 16911 14977
rect 17586 14968 17592 14980
rect 17644 14968 17650 15020
rect 18141 15011 18199 15017
rect 18141 14977 18153 15011
rect 18187 15008 18199 15011
rect 18248 15008 18276 15036
rect 18187 14980 18276 15008
rect 18417 15011 18475 15017
rect 18187 14977 18199 14980
rect 18141 14971 18199 14977
rect 18417 14977 18429 15011
rect 18463 15008 18475 15011
rect 19978 15008 19984 15020
rect 18463 14980 19984 15008
rect 18463 14977 18475 14980
rect 18417 14971 18475 14977
rect 19978 14968 19984 14980
rect 20036 14968 20042 15020
rect 20257 15011 20315 15017
rect 20257 14977 20269 15011
rect 20303 15008 20315 15011
rect 20346 15008 20352 15020
rect 20303 14980 20352 15008
rect 20303 14977 20315 14980
rect 20257 14971 20315 14977
rect 20346 14968 20352 14980
rect 20404 14968 20410 15020
rect 10652 14912 13124 14940
rect 10652 14900 10658 14912
rect 13170 14900 13176 14952
rect 13228 14940 13234 14952
rect 13228 14912 13273 14940
rect 13228 14900 13234 14912
rect 19150 14900 19156 14952
rect 19208 14940 19214 14952
rect 20073 14943 20131 14949
rect 20073 14940 20085 14943
rect 19208 14912 20085 14940
rect 19208 14900 19214 14912
rect 20073 14909 20085 14912
rect 20119 14909 20131 14943
rect 21008 14940 21036 15036
rect 22097 15011 22155 15017
rect 22097 14977 22109 15011
rect 22143 15008 22155 15011
rect 23106 15008 23112 15020
rect 22143 14980 23112 15008
rect 22143 14977 22155 14980
rect 22097 14971 22155 14977
rect 23106 14968 23112 14980
rect 23164 14968 23170 15020
rect 24412 15008 24440 15048
rect 24228 14980 24440 15008
rect 24673 15011 24731 15017
rect 22370 14940 22376 14952
rect 21008 14912 22376 14940
rect 20073 14903 20131 14909
rect 22370 14900 22376 14912
rect 22428 14900 22434 14952
rect 22557 14943 22615 14949
rect 22557 14909 22569 14943
rect 22603 14909 22615 14943
rect 22557 14903 22615 14909
rect 10962 14804 10968 14816
rect 8956 14776 10968 14804
rect 10962 14764 10968 14776
rect 11020 14764 11026 14816
rect 11698 14764 11704 14816
rect 11756 14804 11762 14816
rect 11885 14807 11943 14813
rect 11885 14804 11897 14807
rect 11756 14776 11897 14804
rect 11756 14764 11762 14776
rect 11885 14773 11897 14776
rect 11931 14773 11943 14807
rect 14550 14804 14556 14816
rect 14511 14776 14556 14804
rect 11885 14767 11943 14773
rect 14550 14764 14556 14776
rect 14608 14764 14614 14816
rect 18966 14764 18972 14816
rect 19024 14804 19030 14816
rect 19153 14807 19211 14813
rect 19153 14804 19165 14807
rect 19024 14776 19165 14804
rect 19024 14764 19030 14776
rect 19153 14773 19165 14776
rect 19199 14773 19211 14807
rect 20438 14804 20444 14816
rect 20399 14776 20444 14804
rect 19153 14767 19211 14773
rect 20438 14764 20444 14776
rect 20496 14764 20502 14816
rect 21082 14804 21088 14816
rect 21043 14776 21088 14804
rect 21082 14764 21088 14776
rect 21140 14764 21146 14816
rect 21358 14764 21364 14816
rect 21416 14804 21422 14816
rect 22572 14804 22600 14903
rect 24228 14804 24256 14980
rect 24673 14977 24685 15011
rect 24719 15008 24731 15011
rect 25314 15008 25320 15020
rect 24719 14980 25320 15008
rect 24719 14977 24731 14980
rect 24673 14971 24731 14977
rect 25314 14968 25320 14980
rect 25372 14968 25378 15020
rect 25685 15011 25743 15017
rect 25685 14977 25697 15011
rect 25731 15008 25743 15011
rect 26050 15008 26056 15020
rect 25731 14980 26056 15008
rect 25731 14977 25743 14980
rect 25685 14971 25743 14977
rect 24302 14900 24308 14952
rect 24360 14940 24366 14952
rect 24949 14943 25007 14949
rect 24949 14940 24961 14943
rect 24360 14912 24961 14940
rect 24360 14900 24366 14912
rect 24949 14909 24961 14912
rect 24995 14940 25007 14943
rect 25222 14940 25228 14952
rect 24995 14912 25228 14940
rect 24995 14909 25007 14912
rect 24949 14903 25007 14909
rect 25222 14900 25228 14912
rect 25280 14900 25286 14952
rect 25406 14940 25412 14952
rect 25367 14912 25412 14940
rect 25406 14900 25412 14912
rect 25464 14900 25470 14952
rect 24857 14875 24915 14881
rect 24857 14841 24869 14875
rect 24903 14872 24915 14875
rect 25038 14872 25044 14884
rect 24903 14844 25044 14872
rect 24903 14841 24915 14844
rect 24857 14835 24915 14841
rect 25038 14832 25044 14844
rect 25096 14872 25102 14884
rect 25700 14872 25728 14971
rect 26050 14968 26056 14980
rect 26108 14968 26114 15020
rect 25096 14844 25728 14872
rect 25096 14832 25102 14844
rect 21416 14776 24256 14804
rect 24489 14807 24547 14813
rect 21416 14764 21422 14776
rect 24489 14773 24501 14807
rect 24535 14804 24547 14807
rect 25958 14804 25964 14816
rect 24535 14776 25964 14804
rect 24535 14773 24547 14776
rect 24489 14767 24547 14773
rect 25958 14764 25964 14776
rect 26016 14764 26022 14816
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 7006 14600 7012 14612
rect 6840 14572 7012 14600
rect 6840 14473 6868 14572
rect 7006 14560 7012 14572
rect 7064 14560 7070 14612
rect 9582 14560 9588 14612
rect 9640 14600 9646 14612
rect 9677 14603 9735 14609
rect 9677 14600 9689 14603
rect 9640 14572 9689 14600
rect 9640 14560 9646 14572
rect 9677 14569 9689 14572
rect 9723 14569 9735 14603
rect 9677 14563 9735 14569
rect 9766 14560 9772 14612
rect 9824 14600 9830 14612
rect 9861 14603 9919 14609
rect 9861 14600 9873 14603
rect 9824 14572 9873 14600
rect 9824 14560 9830 14572
rect 9861 14569 9873 14572
rect 9907 14569 9919 14603
rect 10594 14600 10600 14612
rect 10555 14572 10600 14600
rect 9861 14563 9919 14569
rect 10594 14560 10600 14572
rect 10652 14560 10658 14612
rect 10781 14603 10839 14609
rect 10781 14569 10793 14603
rect 10827 14600 10839 14603
rect 10870 14600 10876 14612
rect 10827 14572 10876 14600
rect 10827 14569 10839 14572
rect 10781 14563 10839 14569
rect 10870 14560 10876 14572
rect 10928 14560 10934 14612
rect 13078 14600 13084 14612
rect 13039 14572 13084 14600
rect 13078 14560 13084 14572
rect 13136 14560 13142 14612
rect 15378 14560 15384 14612
rect 15436 14600 15442 14612
rect 16390 14600 16396 14612
rect 15436 14572 16396 14600
rect 15436 14560 15442 14572
rect 16390 14560 16396 14572
rect 16448 14560 16454 14612
rect 18693 14603 18751 14609
rect 18693 14569 18705 14603
rect 18739 14600 18751 14603
rect 18874 14600 18880 14612
rect 18739 14572 18880 14600
rect 18739 14569 18751 14572
rect 18693 14563 18751 14569
rect 18874 14560 18880 14572
rect 18932 14600 18938 14612
rect 23106 14600 23112 14612
rect 18932 14572 22094 14600
rect 23067 14572 23112 14600
rect 18932 14560 18938 14572
rect 22066 14532 22094 14572
rect 23106 14560 23112 14572
rect 23164 14560 23170 14612
rect 23934 14560 23940 14612
rect 23992 14600 23998 14612
rect 23992 14572 24900 14600
rect 23992 14560 23998 14572
rect 22066 14504 24808 14532
rect 6825 14467 6883 14473
rect 6825 14433 6837 14467
rect 6871 14433 6883 14467
rect 6825 14427 6883 14433
rect 9950 14424 9956 14476
rect 10008 14464 10014 14476
rect 10413 14467 10471 14473
rect 10413 14464 10425 14467
rect 10008 14436 10425 14464
rect 10008 14424 10014 14436
rect 10413 14433 10425 14436
rect 10459 14433 10471 14467
rect 10413 14427 10471 14433
rect 11054 14424 11060 14476
rect 11112 14464 11118 14476
rect 14185 14467 14243 14473
rect 11112 14436 11836 14464
rect 11112 14424 11118 14436
rect 6914 14356 6920 14408
rect 6972 14396 6978 14408
rect 7081 14399 7139 14405
rect 7081 14396 7093 14399
rect 6972 14368 7093 14396
rect 6972 14356 6978 14368
rect 7081 14365 7093 14368
rect 7127 14365 7139 14399
rect 10597 14399 10655 14405
rect 10597 14396 10609 14399
rect 7081 14359 7139 14365
rect 9508 14368 10609 14396
rect 9508 14337 9536 14368
rect 10597 14365 10609 14368
rect 10643 14396 10655 14399
rect 10962 14396 10968 14408
rect 10643 14368 10968 14396
rect 10643 14365 10655 14368
rect 10597 14359 10655 14365
rect 10962 14356 10968 14368
rect 11020 14356 11026 14408
rect 11701 14399 11759 14405
rect 11701 14365 11713 14399
rect 11747 14365 11759 14399
rect 11808 14396 11836 14436
rect 14185 14433 14197 14467
rect 14231 14464 14243 14467
rect 14550 14464 14556 14476
rect 14231 14436 14556 14464
rect 14231 14433 14243 14436
rect 14185 14427 14243 14433
rect 14550 14424 14556 14436
rect 14608 14464 14614 14476
rect 22278 14464 22284 14476
rect 14608 14436 15148 14464
rect 14608 14424 14614 14436
rect 11957 14399 12015 14405
rect 11957 14396 11969 14399
rect 11808 14368 11969 14396
rect 11701 14359 11759 14365
rect 11957 14365 11969 14368
rect 12003 14365 12015 14399
rect 11957 14359 12015 14365
rect 9493 14331 9551 14337
rect 9493 14297 9505 14331
rect 9539 14297 9551 14331
rect 9493 14291 9551 14297
rect 9582 14288 9588 14340
rect 9640 14328 9646 14340
rect 10321 14331 10379 14337
rect 10321 14328 10333 14331
rect 9640 14300 10333 14328
rect 9640 14288 9646 14300
rect 10321 14297 10333 14300
rect 10367 14297 10379 14331
rect 10321 14291 10379 14297
rect 11514 14288 11520 14340
rect 11572 14328 11578 14340
rect 11716 14328 11744 14359
rect 12434 14356 12440 14408
rect 12492 14396 12498 14408
rect 12894 14396 12900 14408
rect 12492 14368 12900 14396
rect 12492 14356 12498 14368
rect 12894 14356 12900 14368
rect 12952 14396 12958 14408
rect 15010 14405 15016 14408
rect 14369 14399 14427 14405
rect 14369 14396 14381 14399
rect 12952 14368 14381 14396
rect 12952 14356 12958 14368
rect 14369 14365 14381 14368
rect 14415 14365 14427 14399
rect 15002 14399 15016 14405
rect 15002 14398 15014 14399
rect 14997 14396 15014 14398
rect 14927 14368 15014 14396
rect 14369 14359 14427 14365
rect 14997 14365 15014 14368
rect 14997 14356 15016 14365
rect 15068 14356 15074 14408
rect 15120 14396 15148 14436
rect 22204 14436 22284 14464
rect 15562 14396 15568 14408
rect 15120 14368 15568 14396
rect 15562 14356 15568 14368
rect 15620 14356 15626 14408
rect 17310 14396 17316 14408
rect 17271 14368 17316 14396
rect 17310 14356 17316 14368
rect 17368 14356 17374 14408
rect 19426 14396 19432 14408
rect 19387 14368 19432 14396
rect 19426 14356 19432 14368
rect 19484 14356 19490 14408
rect 20073 14399 20131 14405
rect 20073 14365 20085 14399
rect 20119 14396 20131 14399
rect 21358 14396 21364 14408
rect 20119 14368 21364 14396
rect 20119 14365 20131 14368
rect 20073 14359 20131 14365
rect 21358 14356 21364 14368
rect 21416 14356 21422 14408
rect 21913 14399 21971 14405
rect 21913 14365 21925 14399
rect 21959 14365 21971 14399
rect 21913 14359 21971 14365
rect 22097 14399 22155 14405
rect 22097 14365 22109 14399
rect 22143 14396 22155 14399
rect 22204 14396 22232 14436
rect 22278 14424 22284 14436
rect 22336 14424 22342 14476
rect 22462 14424 22468 14476
rect 22520 14464 22526 14476
rect 22520 14436 22968 14464
rect 22520 14424 22526 14436
rect 22738 14396 22744 14408
rect 22143 14368 22232 14396
rect 22699 14368 22744 14396
rect 22143 14365 22155 14368
rect 22097 14359 22155 14365
rect 13170 14328 13176 14340
rect 11572 14300 13176 14328
rect 11572 14288 11578 14300
rect 13170 14288 13176 14300
rect 13228 14328 13234 14340
rect 14997 14328 15025 14356
rect 15286 14337 15292 14340
rect 13228 14300 15025 14328
rect 13228 14288 13234 14300
rect 15280 14291 15292 14337
rect 15344 14328 15350 14340
rect 17580 14331 17638 14337
rect 15344 14300 15380 14328
rect 15286 14288 15292 14291
rect 15344 14288 15350 14300
rect 17580 14297 17592 14331
rect 17626 14328 17638 14331
rect 17626 14300 19288 14328
rect 17626 14297 17638 14300
rect 17580 14291 17638 14297
rect 8205 14263 8263 14269
rect 8205 14229 8217 14263
rect 8251 14260 8263 14263
rect 8294 14260 8300 14272
rect 8251 14232 8300 14260
rect 8251 14229 8263 14232
rect 8205 14223 8263 14229
rect 8294 14220 8300 14232
rect 8352 14220 8358 14272
rect 9703 14263 9761 14269
rect 9703 14229 9715 14263
rect 9749 14260 9761 14263
rect 9950 14260 9956 14272
rect 9749 14232 9956 14260
rect 9749 14229 9761 14232
rect 9703 14223 9761 14229
rect 9950 14220 9956 14232
rect 10008 14220 10014 14272
rect 14553 14263 14611 14269
rect 14553 14229 14565 14263
rect 14599 14260 14611 14263
rect 16114 14260 16120 14272
rect 14599 14232 16120 14260
rect 14599 14229 14611 14232
rect 14553 14223 14611 14229
rect 16114 14220 16120 14232
rect 16172 14220 16178 14272
rect 19260 14269 19288 14300
rect 19978 14288 19984 14340
rect 20036 14328 20042 14340
rect 20318 14331 20376 14337
rect 20318 14328 20330 14331
rect 20036 14300 20330 14328
rect 20036 14288 20042 14300
rect 20318 14297 20330 14300
rect 20364 14297 20376 14331
rect 21818 14328 21824 14340
rect 20318 14291 20376 14297
rect 21284 14300 21824 14328
rect 19245 14263 19303 14269
rect 19245 14229 19257 14263
rect 19291 14229 19303 14263
rect 19245 14223 19303 14229
rect 19334 14220 19340 14272
rect 19392 14260 19398 14272
rect 21284 14260 21312 14300
rect 21818 14288 21824 14300
rect 21876 14328 21882 14340
rect 21928 14328 21956 14359
rect 22738 14356 22744 14368
rect 22796 14356 22802 14408
rect 22940 14405 22968 14436
rect 22925 14399 22983 14405
rect 22925 14365 22937 14399
rect 22971 14365 22983 14399
rect 22925 14359 22983 14365
rect 23569 14399 23627 14405
rect 23569 14365 23581 14399
rect 23615 14396 23627 14399
rect 24670 14396 24676 14408
rect 23615 14368 24676 14396
rect 23615 14365 23627 14368
rect 23569 14359 23627 14365
rect 24670 14356 24676 14368
rect 24728 14356 24734 14408
rect 24780 14405 24808 14504
rect 24872 14473 24900 14572
rect 24857 14467 24915 14473
rect 24857 14433 24869 14467
rect 24903 14433 24915 14467
rect 25038 14464 25044 14476
rect 24999 14436 25044 14464
rect 24857 14427 24915 14433
rect 25038 14424 25044 14436
rect 25096 14424 25102 14476
rect 25682 14424 25688 14476
rect 25740 14464 25746 14476
rect 25961 14467 26019 14473
rect 25961 14464 25973 14467
rect 25740 14436 25973 14464
rect 25740 14424 25746 14436
rect 25961 14433 25973 14436
rect 26007 14433 26019 14467
rect 25961 14427 26019 14433
rect 26234 14405 26240 14408
rect 24765 14399 24823 14405
rect 24765 14365 24777 14399
rect 24811 14365 24823 14399
rect 26228 14396 26240 14405
rect 26195 14368 26240 14396
rect 24765 14359 24823 14365
rect 26228 14359 26240 14368
rect 26234 14356 26240 14359
rect 26292 14356 26298 14408
rect 24302 14328 24308 14340
rect 21876 14300 21956 14328
rect 22066 14300 24308 14328
rect 21876 14288 21882 14300
rect 21450 14260 21456 14272
rect 19392 14232 21312 14260
rect 21411 14232 21456 14260
rect 19392 14220 19398 14232
rect 21450 14220 21456 14232
rect 21508 14260 21514 14272
rect 22066 14260 22094 14300
rect 24302 14288 24308 14300
rect 24360 14288 24366 14340
rect 25222 14328 25228 14340
rect 24412 14300 25228 14328
rect 22278 14260 22284 14272
rect 21508 14232 22094 14260
rect 22239 14232 22284 14260
rect 21508 14220 21514 14232
rect 22278 14220 22284 14232
rect 22336 14220 22342 14272
rect 23753 14263 23811 14269
rect 23753 14229 23765 14263
rect 23799 14260 23811 14263
rect 24118 14260 24124 14272
rect 23799 14232 24124 14260
rect 23799 14229 23811 14232
rect 23753 14223 23811 14229
rect 24118 14220 24124 14232
rect 24176 14220 24182 14272
rect 24412 14269 24440 14300
rect 25222 14288 25228 14300
rect 25280 14288 25286 14340
rect 24397 14263 24455 14269
rect 24397 14229 24409 14263
rect 24443 14229 24455 14263
rect 24397 14223 24455 14229
rect 25406 14220 25412 14272
rect 25464 14260 25470 14272
rect 27341 14263 27399 14269
rect 27341 14260 27353 14263
rect 25464 14232 27353 14260
rect 25464 14220 25470 14232
rect 27341 14229 27353 14232
rect 27387 14260 27399 14263
rect 37734 14260 37740 14272
rect 27387 14232 37740 14260
rect 27387 14229 27399 14232
rect 27341 14223 27399 14229
rect 37734 14220 37740 14232
rect 37792 14220 37798 14272
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 9950 14056 9956 14068
rect 9911 14028 9956 14056
rect 9950 14016 9956 14028
rect 10008 14016 10014 14068
rect 10226 14016 10232 14068
rect 10284 14056 10290 14068
rect 11517 14059 11575 14065
rect 11517 14056 11529 14059
rect 10284 14028 11529 14056
rect 10284 14016 10290 14028
rect 11517 14025 11529 14028
rect 11563 14025 11575 14059
rect 11517 14019 11575 14025
rect 12710 14016 12716 14068
rect 12768 14056 12774 14068
rect 13633 14059 13691 14065
rect 13633 14056 13645 14059
rect 12768 14028 13645 14056
rect 12768 14016 12774 14028
rect 13633 14025 13645 14028
rect 13679 14025 13691 14059
rect 18966 14056 18972 14068
rect 13633 14019 13691 14025
rect 15028 14028 15516 14056
rect 18927 14028 18972 14056
rect 8294 13988 8300 14000
rect 7944 13960 8300 13988
rect 7944 13929 7972 13960
rect 8294 13948 8300 13960
rect 8352 13988 8358 14000
rect 9766 13988 9772 14000
rect 8352 13960 9628 13988
rect 9727 13960 9772 13988
rect 8352 13948 8358 13960
rect 9600 13932 9628 13960
rect 9766 13948 9772 13960
rect 9824 13948 9830 14000
rect 11606 13988 11612 14000
rect 10612 13960 11612 13988
rect 7929 13923 7987 13929
rect 7929 13889 7941 13923
rect 7975 13889 7987 13923
rect 7929 13883 7987 13889
rect 8018 13880 8024 13932
rect 8076 13920 8082 13932
rect 8754 13920 8760 13932
rect 8076 13892 8616 13920
rect 8715 13892 8760 13920
rect 8076 13880 8082 13892
rect 7745 13855 7803 13861
rect 7745 13821 7757 13855
rect 7791 13852 7803 13855
rect 8036 13852 8064 13880
rect 7791 13824 8064 13852
rect 8113 13855 8171 13861
rect 7791 13821 7803 13824
rect 7745 13815 7803 13821
rect 8113 13821 8125 13855
rect 8159 13852 8171 13855
rect 8478 13852 8484 13864
rect 8159 13824 8484 13852
rect 8159 13821 8171 13824
rect 8113 13815 8171 13821
rect 8478 13812 8484 13824
rect 8536 13812 8542 13864
rect 8588 13861 8616 13892
rect 8754 13880 8760 13892
rect 8812 13920 8818 13932
rect 9401 13923 9459 13929
rect 9401 13920 9413 13923
rect 8812 13892 9413 13920
rect 8812 13880 8818 13892
rect 9401 13889 9413 13892
rect 9447 13889 9459 13923
rect 9582 13920 9588 13932
rect 9543 13892 9588 13920
rect 9401 13883 9459 13889
rect 9582 13880 9588 13892
rect 9640 13880 9646 13932
rect 9674 13880 9680 13932
rect 9732 13920 9738 13932
rect 10612 13929 10640 13960
rect 11606 13948 11612 13960
rect 11664 13988 11670 14000
rect 12437 13991 12495 13997
rect 12437 13988 12449 13991
rect 11664 13960 12449 13988
rect 11664 13948 11670 13960
rect 12437 13957 12449 13960
rect 12483 13988 12495 13991
rect 15028 13988 15056 14028
rect 12483 13960 15056 13988
rect 12483 13957 12495 13960
rect 12437 13951 12495 13957
rect 15378 13948 15384 14000
rect 15436 13948 15442 14000
rect 10597 13923 10655 13929
rect 9732 13892 9777 13920
rect 9732 13880 9738 13892
rect 10597 13889 10609 13923
rect 10643 13889 10655 13923
rect 11698 13920 11704 13932
rect 11659 13892 11704 13920
rect 10597 13883 10655 13889
rect 11698 13880 11704 13892
rect 11756 13880 11762 13932
rect 12253 13923 12311 13929
rect 12253 13889 12265 13923
rect 12299 13920 12311 13923
rect 12618 13920 12624 13932
rect 12299 13892 12624 13920
rect 12299 13889 12311 13892
rect 12253 13883 12311 13889
rect 12618 13880 12624 13892
rect 12676 13920 12682 13932
rect 12894 13920 12900 13932
rect 12676 13892 12900 13920
rect 12676 13880 12682 13892
rect 12894 13880 12900 13892
rect 12952 13880 12958 13932
rect 13446 13920 13452 13932
rect 13407 13892 13452 13920
rect 13446 13880 13452 13892
rect 13504 13880 13510 13932
rect 15102 13920 15108 13932
rect 15063 13892 15108 13920
rect 15102 13880 15108 13892
rect 15160 13880 15166 13932
rect 15197 13923 15255 13929
rect 15197 13889 15209 13923
rect 15243 13889 15255 13923
rect 15197 13883 15255 13889
rect 15289 13923 15347 13929
rect 15289 13889 15301 13923
rect 15335 13920 15347 13923
rect 15396 13920 15424 13948
rect 15488 13929 15516 14028
rect 18966 14016 18972 14028
rect 19024 14016 19030 14068
rect 19705 14059 19763 14065
rect 19705 14025 19717 14059
rect 19751 14056 19763 14059
rect 19978 14056 19984 14068
rect 19751 14028 19984 14056
rect 19751 14025 19763 14028
rect 19705 14019 19763 14025
rect 19978 14016 19984 14028
rect 20036 14016 20042 14068
rect 20346 14056 20352 14068
rect 20307 14028 20352 14056
rect 20346 14016 20352 14028
rect 20404 14016 20410 14068
rect 20717 14059 20775 14065
rect 20717 14025 20729 14059
rect 20763 14056 20775 14059
rect 21450 14056 21456 14068
rect 20763 14028 21456 14056
rect 20763 14025 20775 14028
rect 20717 14019 20775 14025
rect 21450 14016 21456 14028
rect 21508 14016 21514 14068
rect 22005 14059 22063 14065
rect 22005 14025 22017 14059
rect 22051 14056 22063 14059
rect 22186 14056 22192 14068
rect 22051 14028 22192 14056
rect 22051 14025 22063 14028
rect 22005 14019 22063 14025
rect 22186 14016 22192 14028
rect 22244 14016 22250 14068
rect 22465 14059 22523 14065
rect 22465 14025 22477 14059
rect 22511 14056 22523 14059
rect 22830 14056 22836 14068
rect 22511 14028 22836 14056
rect 22511 14025 22523 14028
rect 22465 14019 22523 14025
rect 22830 14016 22836 14028
rect 22888 14016 22894 14068
rect 25409 14059 25467 14065
rect 25409 14025 25421 14059
rect 25455 14056 25467 14059
rect 26510 14056 26516 14068
rect 25455 14028 26516 14056
rect 25455 14025 25467 14028
rect 25409 14019 25467 14025
rect 26510 14016 26516 14028
rect 26568 14016 26574 14068
rect 18874 13988 18880 14000
rect 18835 13960 18880 13988
rect 18874 13948 18880 13960
rect 18932 13948 18938 14000
rect 20806 13988 20812 14000
rect 20767 13960 20812 13988
rect 20806 13948 20812 13960
rect 20864 13948 20870 14000
rect 24854 13948 24860 14000
rect 24912 13988 24918 14000
rect 25225 13991 25283 13997
rect 25225 13988 25237 13991
rect 24912 13960 25237 13988
rect 24912 13948 24918 13960
rect 25225 13957 25237 13960
rect 25271 13988 25283 13991
rect 25498 13988 25504 14000
rect 25271 13960 25504 13988
rect 25271 13957 25283 13960
rect 25225 13951 25283 13957
rect 25498 13948 25504 13960
rect 25556 13948 25562 14000
rect 25869 13991 25927 13997
rect 25869 13957 25881 13991
rect 25915 13957 25927 13991
rect 25869 13951 25927 13957
rect 15335 13892 15424 13920
rect 15473 13923 15531 13929
rect 15335 13889 15347 13892
rect 15289 13883 15347 13889
rect 15473 13889 15485 13923
rect 15519 13889 15531 13923
rect 16114 13920 16120 13932
rect 16075 13892 16120 13920
rect 15473 13883 15531 13889
rect 8573 13855 8631 13861
rect 8573 13821 8585 13855
rect 8619 13852 8631 13855
rect 8941 13855 8999 13861
rect 8619 13824 8892 13852
rect 8619 13821 8631 13824
rect 8573 13815 8631 13821
rect 8864 13784 8892 13824
rect 8941 13821 8953 13855
rect 8987 13852 8999 13855
rect 9122 13852 9128 13864
rect 8987 13824 9128 13852
rect 8987 13821 8999 13824
rect 8941 13815 8999 13821
rect 9122 13812 9128 13824
rect 9180 13812 9186 13864
rect 13262 13852 13268 13864
rect 9232 13824 10456 13852
rect 13223 13824 13268 13852
rect 9232 13784 9260 13824
rect 10428 13793 10456 13824
rect 13262 13812 13268 13824
rect 13320 13812 13326 13864
rect 15212 13852 15240 13883
rect 15378 13852 15384 13864
rect 15212 13824 15384 13852
rect 15378 13812 15384 13824
rect 15436 13812 15442 13864
rect 15488 13852 15516 13883
rect 16114 13880 16120 13892
rect 16172 13880 16178 13932
rect 17037 13923 17095 13929
rect 17037 13889 17049 13923
rect 17083 13920 17095 13923
rect 17126 13920 17132 13932
rect 17083 13892 17132 13920
rect 17083 13889 17095 13892
rect 17037 13883 17095 13889
rect 17052 13852 17080 13883
rect 17126 13880 17132 13892
rect 17184 13880 17190 13932
rect 17313 13923 17371 13929
rect 17313 13889 17325 13923
rect 17359 13920 17371 13923
rect 18046 13920 18052 13932
rect 17359 13892 18052 13920
rect 17359 13889 17371 13892
rect 17313 13883 17371 13889
rect 18046 13880 18052 13892
rect 18104 13880 18110 13932
rect 19889 13923 19947 13929
rect 19889 13889 19901 13923
rect 19935 13920 19947 13923
rect 20438 13920 20444 13932
rect 19935 13892 20444 13920
rect 19935 13889 19947 13892
rect 19889 13883 19947 13889
rect 20438 13880 20444 13892
rect 20496 13880 20502 13932
rect 22370 13920 22376 13932
rect 22331 13892 22376 13920
rect 22370 13880 22376 13892
rect 22428 13880 22434 13932
rect 24118 13920 24124 13932
rect 24079 13892 24124 13920
rect 24118 13880 24124 13892
rect 24176 13920 24182 13932
rect 24946 13920 24952 13932
rect 24176 13892 24952 13920
rect 24176 13880 24182 13892
rect 24946 13880 24952 13892
rect 25004 13880 25010 13932
rect 25038 13880 25044 13932
rect 25096 13920 25102 13932
rect 25884 13920 25912 13951
rect 26050 13948 26056 14000
rect 26108 13997 26114 14000
rect 26108 13991 26127 13997
rect 26115 13957 26127 13991
rect 28169 13991 28227 13997
rect 28169 13988 28181 13991
rect 26108 13951 26127 13957
rect 26160 13960 28181 13988
rect 26108 13948 26114 13951
rect 26160 13920 26188 13960
rect 28169 13957 28181 13960
rect 28215 13957 28227 13991
rect 28169 13951 28227 13957
rect 25096 13892 26188 13920
rect 27433 13923 27491 13929
rect 25096 13880 25102 13892
rect 27433 13889 27445 13923
rect 27479 13920 27491 13923
rect 28077 13923 28135 13929
rect 28077 13920 28089 13923
rect 27479 13892 28089 13920
rect 27479 13889 27491 13892
rect 27433 13883 27491 13889
rect 28077 13889 28089 13892
rect 28123 13889 28135 13923
rect 28077 13883 28135 13889
rect 15488 13824 17080 13852
rect 19061 13855 19119 13861
rect 19061 13821 19073 13855
rect 19107 13821 19119 13855
rect 19061 13815 19119 13821
rect 20901 13855 20959 13861
rect 20901 13821 20913 13855
rect 20947 13852 20959 13855
rect 21082 13852 21088 13864
rect 20947 13824 21088 13852
rect 20947 13821 20959 13824
rect 20901 13815 20959 13821
rect 8864 13756 9260 13784
rect 10413 13787 10471 13793
rect 10413 13753 10425 13787
rect 10459 13753 10471 13787
rect 10413 13747 10471 13753
rect 11790 13744 11796 13796
rect 11848 13784 11854 13796
rect 17954 13784 17960 13796
rect 11848 13756 15164 13784
rect 11848 13744 11854 13756
rect 3786 13676 3792 13728
rect 3844 13716 3850 13728
rect 10226 13716 10232 13728
rect 3844 13688 10232 13716
rect 3844 13676 3850 13688
rect 10226 13676 10232 13688
rect 10284 13676 10290 13728
rect 14829 13719 14887 13725
rect 14829 13685 14841 13719
rect 14875 13716 14887 13719
rect 14918 13716 14924 13728
rect 14875 13688 14924 13716
rect 14875 13685 14887 13688
rect 14829 13679 14887 13685
rect 14918 13676 14924 13688
rect 14976 13676 14982 13728
rect 15136 13716 15164 13756
rect 15672 13756 17960 13784
rect 15672 13716 15700 13756
rect 17954 13744 17960 13756
rect 18012 13744 18018 13796
rect 18598 13744 18604 13796
rect 18656 13784 18662 13796
rect 19076 13784 19104 13815
rect 20916 13784 20944 13815
rect 21082 13812 21088 13824
rect 21140 13812 21146 13864
rect 22462 13812 22468 13864
rect 22520 13852 22526 13864
rect 22557 13855 22615 13861
rect 22557 13852 22569 13855
rect 22520 13824 22569 13852
rect 22520 13812 22526 13824
rect 22557 13821 22569 13824
rect 22603 13821 22615 13855
rect 23750 13852 23756 13864
rect 23711 13824 23756 13852
rect 22557 13815 22615 13821
rect 23750 13812 23756 13824
rect 23808 13812 23814 13864
rect 24210 13812 24216 13864
rect 24268 13852 24274 13864
rect 24857 13855 24915 13861
rect 24268 13824 24313 13852
rect 24268 13812 24274 13824
rect 24857 13821 24869 13855
rect 24903 13852 24915 13855
rect 24903 13824 25176 13852
rect 24903 13821 24915 13824
rect 24857 13815 24915 13821
rect 18656 13756 20944 13784
rect 25148 13784 25176 13824
rect 25222 13812 25228 13864
rect 25280 13852 25286 13864
rect 27448 13852 27476 13883
rect 25280 13824 27476 13852
rect 25280 13812 25286 13824
rect 26786 13784 26792 13796
rect 25148 13756 26792 13784
rect 18656 13744 18662 13756
rect 26786 13744 26792 13756
rect 26844 13744 26850 13796
rect 27614 13784 27620 13796
rect 27575 13756 27620 13784
rect 27614 13744 27620 13756
rect 27672 13744 27678 13796
rect 15136 13688 15700 13716
rect 15746 13676 15752 13728
rect 15804 13716 15810 13728
rect 15933 13719 15991 13725
rect 15933 13716 15945 13719
rect 15804 13688 15945 13716
rect 15804 13676 15810 13688
rect 15933 13685 15945 13688
rect 15979 13685 15991 13719
rect 15933 13679 15991 13685
rect 18046 13676 18052 13728
rect 18104 13716 18110 13728
rect 18509 13719 18567 13725
rect 18509 13716 18521 13719
rect 18104 13688 18521 13716
rect 18104 13676 18110 13688
rect 18509 13685 18521 13688
rect 18555 13685 18567 13719
rect 18509 13679 18567 13685
rect 23658 13676 23664 13728
rect 23716 13716 23722 13728
rect 24397 13719 24455 13725
rect 24397 13716 24409 13719
rect 23716 13688 24409 13716
rect 23716 13676 23722 13688
rect 24397 13685 24409 13688
rect 24443 13685 24455 13719
rect 25222 13716 25228 13728
rect 25183 13688 25228 13716
rect 24397 13679 24455 13685
rect 25222 13676 25228 13688
rect 25280 13676 25286 13728
rect 25958 13676 25964 13728
rect 26016 13716 26022 13728
rect 26053 13719 26111 13725
rect 26053 13716 26065 13719
rect 26016 13688 26065 13716
rect 26016 13676 26022 13688
rect 26053 13685 26065 13688
rect 26099 13716 26111 13719
rect 26142 13716 26148 13728
rect 26099 13688 26148 13716
rect 26099 13685 26111 13688
rect 26053 13679 26111 13685
rect 26142 13676 26148 13688
rect 26200 13676 26206 13728
rect 26237 13719 26295 13725
rect 26237 13685 26249 13719
rect 26283 13716 26295 13719
rect 26418 13716 26424 13728
rect 26283 13688 26424 13716
rect 26283 13685 26295 13688
rect 26237 13679 26295 13685
rect 26418 13676 26424 13688
rect 26476 13676 26482 13728
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 8389 13515 8447 13521
rect 8389 13481 8401 13515
rect 8435 13512 8447 13515
rect 8754 13512 8760 13524
rect 8435 13484 8760 13512
rect 8435 13481 8447 13484
rect 8389 13475 8447 13481
rect 8754 13472 8760 13484
rect 8812 13472 8818 13524
rect 9582 13472 9588 13524
rect 9640 13512 9646 13524
rect 9677 13515 9735 13521
rect 9677 13512 9689 13515
rect 9640 13484 9689 13512
rect 9640 13472 9646 13484
rect 9677 13481 9689 13484
rect 9723 13481 9735 13515
rect 10134 13512 10140 13524
rect 10095 13484 10140 13512
rect 9677 13475 9735 13481
rect 10134 13472 10140 13484
rect 10192 13472 10198 13524
rect 10226 13472 10232 13524
rect 10284 13512 10290 13524
rect 10284 13484 26556 13512
rect 10284 13472 10290 13484
rect 8772 13444 8800 13472
rect 14461 13447 14519 13453
rect 8772 13416 9996 13444
rect 7006 13376 7012 13388
rect 6967 13348 7012 13376
rect 7006 13336 7012 13348
rect 7064 13336 7070 13388
rect 9674 13336 9680 13388
rect 9732 13376 9738 13388
rect 9769 13379 9827 13385
rect 9769 13376 9781 13379
rect 9732 13348 9781 13376
rect 9732 13336 9738 13348
rect 9769 13345 9781 13348
rect 9815 13345 9827 13379
rect 9769 13339 9827 13345
rect 8478 13268 8484 13320
rect 8536 13308 8542 13320
rect 9968 13317 9996 13416
rect 14461 13413 14473 13447
rect 14507 13444 14519 13447
rect 15286 13444 15292 13456
rect 14507 13416 15292 13444
rect 14507 13413 14519 13416
rect 14461 13407 14519 13413
rect 15286 13404 15292 13416
rect 15344 13404 15350 13456
rect 18233 13447 18291 13453
rect 18233 13413 18245 13447
rect 18279 13444 18291 13447
rect 19426 13444 19432 13456
rect 18279 13416 19432 13444
rect 18279 13413 18291 13416
rect 18233 13407 18291 13413
rect 19426 13404 19432 13416
rect 19484 13404 19490 13456
rect 24946 13404 24952 13456
rect 25004 13444 25010 13456
rect 25590 13444 25596 13456
rect 25004 13416 25596 13444
rect 25004 13404 25010 13416
rect 25590 13404 25596 13416
rect 25648 13444 25654 13456
rect 26142 13444 26148 13456
rect 25648 13416 26148 13444
rect 25648 13404 25654 13416
rect 26142 13404 26148 13416
rect 26200 13404 26206 13456
rect 26528 13453 26556 13484
rect 26513 13447 26571 13453
rect 26513 13413 26525 13447
rect 26559 13413 26571 13447
rect 26513 13407 26571 13413
rect 13541 13379 13599 13385
rect 13541 13376 13553 13379
rect 12728 13348 13553 13376
rect 9125 13311 9183 13317
rect 9125 13308 9137 13311
rect 8536 13280 9137 13308
rect 8536 13268 8542 13280
rect 9125 13277 9137 13280
rect 9171 13277 9183 13311
rect 9125 13271 9183 13277
rect 9953 13311 10011 13317
rect 9953 13277 9965 13311
rect 9999 13277 10011 13311
rect 11606 13308 11612 13320
rect 11567 13280 11612 13308
rect 9953 13271 10011 13277
rect 11606 13268 11612 13280
rect 11664 13268 11670 13320
rect 12728 13317 12756 13348
rect 13541 13345 13553 13348
rect 13587 13345 13599 13379
rect 13541 13339 13599 13345
rect 14550 13336 14556 13388
rect 14608 13376 14614 13388
rect 14829 13379 14887 13385
rect 14829 13376 14841 13379
rect 14608 13348 14841 13376
rect 14608 13336 14614 13348
rect 14829 13345 14841 13348
rect 14875 13345 14887 13379
rect 14829 13339 14887 13345
rect 15102 13336 15108 13388
rect 15160 13376 15166 13388
rect 15473 13379 15531 13385
rect 15473 13376 15485 13379
rect 15160 13348 15485 13376
rect 15160 13336 15166 13348
rect 15473 13345 15485 13348
rect 15519 13345 15531 13379
rect 15473 13339 15531 13345
rect 17865 13379 17923 13385
rect 17865 13345 17877 13379
rect 17911 13376 17923 13379
rect 17954 13376 17960 13388
rect 17911 13348 17960 13376
rect 17911 13345 17923 13348
rect 17865 13339 17923 13345
rect 17954 13336 17960 13348
rect 18012 13336 18018 13388
rect 18138 13336 18144 13388
rect 18196 13376 18202 13388
rect 19242 13376 19248 13388
rect 18196 13348 19248 13376
rect 18196 13336 18202 13348
rect 19242 13336 19248 13348
rect 19300 13336 19306 13388
rect 25038 13376 25044 13388
rect 21008 13348 21588 13376
rect 12713 13311 12771 13317
rect 12713 13277 12725 13311
rect 12759 13277 12771 13311
rect 12713 13271 12771 13277
rect 13265 13311 13323 13317
rect 13265 13277 13277 13311
rect 13311 13277 13323 13311
rect 13265 13271 13323 13277
rect 13357 13311 13415 13317
rect 13357 13277 13369 13311
rect 13403 13308 13415 13311
rect 13446 13308 13452 13320
rect 13403 13280 13452 13308
rect 13403 13277 13415 13280
rect 13357 13271 13415 13277
rect 7276 13243 7334 13249
rect 7276 13209 7288 13243
rect 7322 13240 7334 13243
rect 9677 13243 9735 13249
rect 7322 13212 8984 13240
rect 7322 13209 7334 13212
rect 7276 13203 7334 13209
rect 8956 13181 8984 13212
rect 9677 13209 9689 13243
rect 9723 13240 9735 13243
rect 9766 13240 9772 13252
rect 9723 13212 9772 13240
rect 9723 13209 9735 13212
rect 9677 13203 9735 13209
rect 9766 13200 9772 13212
rect 9824 13240 9830 13252
rect 10962 13240 10968 13252
rect 9824 13212 10968 13240
rect 9824 13200 9830 13212
rect 10962 13200 10968 13212
rect 11020 13200 11026 13252
rect 11790 13240 11796 13252
rect 11751 13212 11796 13240
rect 11790 13200 11796 13212
rect 11848 13200 11854 13252
rect 13280 13240 13308 13271
rect 13446 13268 13452 13280
rect 13504 13268 13510 13320
rect 14645 13311 14703 13317
rect 14645 13277 14657 13311
rect 14691 13277 14703 13311
rect 14645 13271 14703 13277
rect 14550 13240 14556 13252
rect 13280 13212 14556 13240
rect 14550 13200 14556 13212
rect 14608 13200 14614 13252
rect 8941 13175 8999 13181
rect 8941 13141 8953 13175
rect 8987 13141 8999 13175
rect 12526 13172 12532 13184
rect 12487 13144 12532 13172
rect 8941 13135 8999 13141
rect 12526 13132 12532 13144
rect 12584 13132 12590 13184
rect 14660 13172 14688 13271
rect 14734 13268 14740 13320
rect 14792 13308 14798 13320
rect 14918 13317 14924 13320
rect 14914 13308 14924 13317
rect 14792 13280 14837 13308
rect 14879 13280 14924 13308
rect 14792 13268 14798 13280
rect 14914 13271 14924 13280
rect 14918 13268 14924 13271
rect 14976 13268 14982 13320
rect 15746 13317 15752 13320
rect 15740 13308 15752 13317
rect 15707 13280 15752 13308
rect 15740 13271 15752 13280
rect 15746 13268 15752 13271
rect 15804 13268 15810 13320
rect 18046 13308 18052 13320
rect 18007 13280 18052 13308
rect 18046 13268 18052 13280
rect 18104 13268 18110 13320
rect 19426 13308 19432 13320
rect 19387 13280 19432 13308
rect 19426 13268 19432 13280
rect 19484 13268 19490 13320
rect 21008 13317 21036 13348
rect 20993 13311 21051 13317
rect 20993 13277 21005 13311
rect 21039 13277 21051 13311
rect 20993 13271 21051 13277
rect 21082 13268 21088 13320
rect 21140 13308 21146 13320
rect 21358 13308 21364 13320
rect 21140 13280 21364 13308
rect 21140 13268 21146 13280
rect 21358 13268 21364 13280
rect 21416 13308 21422 13320
rect 21453 13311 21511 13317
rect 21453 13308 21465 13311
rect 21416 13280 21465 13308
rect 21416 13268 21422 13280
rect 21453 13277 21465 13280
rect 21499 13277 21511 13311
rect 21560 13308 21588 13348
rect 23676 13348 25044 13376
rect 22278 13308 22284 13320
rect 21560 13280 22284 13308
rect 21453 13271 21511 13277
rect 22278 13268 22284 13280
rect 22336 13268 22342 13320
rect 23676 13317 23704 13348
rect 25038 13336 25044 13348
rect 25096 13336 25102 13388
rect 25777 13379 25835 13385
rect 25777 13345 25789 13379
rect 25823 13376 25835 13379
rect 25823 13348 26004 13376
rect 25823 13345 25835 13348
rect 25777 13339 25835 13345
rect 23661 13311 23719 13317
rect 23661 13277 23673 13311
rect 23707 13277 23719 13311
rect 23661 13271 23719 13277
rect 24762 13268 24768 13320
rect 24820 13308 24826 13320
rect 24857 13311 24915 13317
rect 24857 13308 24869 13311
rect 24820 13280 24869 13308
rect 24820 13268 24826 13280
rect 24857 13277 24869 13280
rect 24903 13277 24915 13311
rect 24857 13271 24915 13277
rect 25869 13311 25927 13317
rect 25869 13277 25881 13311
rect 25915 13277 25927 13311
rect 25976 13308 26004 13348
rect 26326 13336 26332 13388
rect 26384 13376 26390 13388
rect 27249 13379 27307 13385
rect 27249 13376 27261 13379
rect 26384 13348 27261 13376
rect 26384 13336 26390 13348
rect 27249 13345 27261 13348
rect 27295 13345 27307 13379
rect 27249 13339 27307 13345
rect 25976 13280 26924 13308
rect 25869 13271 25927 13277
rect 16942 13200 16948 13252
rect 17000 13240 17006 13252
rect 19613 13243 19671 13249
rect 19613 13240 19625 13243
rect 17000 13212 19625 13240
rect 17000 13200 17006 13212
rect 19613 13209 19625 13212
rect 19659 13209 19671 13243
rect 21698 13243 21756 13249
rect 21698 13240 21710 13243
rect 19613 13203 19671 13209
rect 20824 13212 21710 13240
rect 15102 13172 15108 13184
rect 14660 13144 15108 13172
rect 15102 13132 15108 13144
rect 15160 13132 15166 13184
rect 15654 13132 15660 13184
rect 15712 13172 15718 13184
rect 16853 13175 16911 13181
rect 16853 13172 16865 13175
rect 15712 13144 16865 13172
rect 15712 13132 15718 13144
rect 16853 13141 16865 13144
rect 16899 13141 16911 13175
rect 16853 13135 16911 13141
rect 17954 13132 17960 13184
rect 18012 13172 18018 13184
rect 19242 13172 19248 13184
rect 18012 13144 19248 13172
rect 18012 13132 18018 13144
rect 19242 13132 19248 13144
rect 19300 13132 19306 13184
rect 20824 13181 20852 13212
rect 21698 13209 21710 13212
rect 21744 13209 21756 13243
rect 21698 13203 21756 13209
rect 23845 13243 23903 13249
rect 23845 13209 23857 13243
rect 23891 13240 23903 13243
rect 25682 13240 25688 13252
rect 23891 13212 25688 13240
rect 23891 13209 23903 13212
rect 23845 13203 23903 13209
rect 25682 13200 25688 13212
rect 25740 13240 25746 13252
rect 25884 13240 25912 13271
rect 25740 13212 25912 13240
rect 25961 13243 26019 13249
rect 25740 13200 25746 13212
rect 25961 13209 25973 13243
rect 26007 13240 26019 13243
rect 26142 13240 26148 13252
rect 26007 13212 26148 13240
rect 26007 13209 26019 13212
rect 25961 13203 26019 13209
rect 26142 13200 26148 13212
rect 26200 13200 26206 13252
rect 26326 13240 26332 13252
rect 26287 13212 26332 13240
rect 26326 13200 26332 13212
rect 26384 13200 26390 13252
rect 26896 13240 26924 13280
rect 26970 13268 26976 13320
rect 27028 13308 27034 13320
rect 27525 13311 27583 13317
rect 27525 13308 27537 13311
rect 27028 13280 27537 13308
rect 27028 13268 27034 13280
rect 27525 13277 27537 13280
rect 27571 13277 27583 13311
rect 27525 13271 27583 13277
rect 27154 13240 27160 13252
rect 26896 13212 27160 13240
rect 27154 13200 27160 13212
rect 27212 13200 27218 13252
rect 20809 13175 20867 13181
rect 20809 13141 20821 13175
rect 20855 13141 20867 13175
rect 20809 13135 20867 13141
rect 22370 13132 22376 13184
rect 22428 13172 22434 13184
rect 22833 13175 22891 13181
rect 22833 13172 22845 13175
rect 22428 13144 22845 13172
rect 22428 13132 22434 13144
rect 22833 13141 22845 13144
rect 22879 13172 22891 13175
rect 23382 13172 23388 13184
rect 22879 13144 23388 13172
rect 22879 13141 22891 13144
rect 22833 13135 22891 13141
rect 23382 13132 23388 13144
rect 23440 13132 23446 13184
rect 24118 13132 24124 13184
rect 24176 13172 24182 13184
rect 24397 13175 24455 13181
rect 24397 13172 24409 13175
rect 24176 13144 24409 13172
rect 24176 13132 24182 13144
rect 24397 13141 24409 13144
rect 24443 13141 24455 13175
rect 24397 13135 24455 13141
rect 24765 13175 24823 13181
rect 24765 13141 24777 13175
rect 24811 13172 24823 13175
rect 24946 13172 24952 13184
rect 24811 13144 24952 13172
rect 24811 13141 24823 13144
rect 24765 13135 24823 13141
rect 24946 13132 24952 13144
rect 25004 13172 25010 13184
rect 25498 13172 25504 13184
rect 25004 13144 25504 13172
rect 25004 13132 25010 13144
rect 25498 13132 25504 13144
rect 25556 13132 25562 13184
rect 25774 13132 25780 13184
rect 25832 13172 25838 13184
rect 27614 13172 27620 13184
rect 25832 13144 27620 13172
rect 25832 13132 25838 13144
rect 27614 13132 27620 13144
rect 27672 13132 27678 13184
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 2746 12940 14504 12968
rect 1486 12860 1492 12912
rect 1544 12900 1550 12912
rect 2746 12900 2774 12940
rect 1544 12872 2774 12900
rect 1544 12860 1550 12872
rect 12526 12860 12532 12912
rect 12584 12900 12590 12912
rect 13602 12903 13660 12909
rect 13602 12900 13614 12903
rect 12584 12872 13614 12900
rect 12584 12860 12590 12872
rect 13602 12869 13614 12872
rect 13648 12869 13660 12903
rect 14476 12900 14504 12940
rect 15470 12928 15476 12980
rect 15528 12968 15534 12980
rect 15657 12971 15715 12977
rect 15657 12968 15669 12971
rect 15528 12940 15669 12968
rect 15528 12928 15534 12940
rect 15657 12937 15669 12940
rect 15703 12937 15715 12971
rect 15657 12931 15715 12937
rect 16669 12971 16727 12977
rect 16669 12937 16681 12971
rect 16715 12937 16727 12971
rect 16669 12931 16727 12937
rect 20073 12971 20131 12977
rect 20073 12937 20085 12971
rect 20119 12968 20131 12971
rect 20254 12968 20260 12980
rect 20119 12940 20260 12968
rect 20119 12937 20131 12940
rect 20073 12931 20131 12937
rect 16684 12900 16712 12931
rect 20254 12928 20260 12940
rect 20312 12928 20318 12980
rect 22094 12928 22100 12980
rect 22152 12968 22158 12980
rect 22281 12971 22339 12977
rect 22281 12968 22293 12971
rect 22152 12940 22293 12968
rect 22152 12928 22158 12940
rect 22281 12937 22293 12940
rect 22327 12937 22339 12971
rect 22281 12931 22339 12937
rect 25777 12971 25835 12977
rect 25777 12937 25789 12971
rect 25823 12968 25835 12971
rect 26326 12968 26332 12980
rect 25823 12940 26332 12968
rect 25823 12937 25835 12940
rect 25777 12931 25835 12937
rect 26326 12928 26332 12940
rect 26384 12928 26390 12980
rect 17558 12903 17616 12909
rect 17558 12900 17570 12903
rect 14476 12872 15783 12900
rect 16684 12872 17570 12900
rect 13602 12863 13660 12869
rect 7006 12792 7012 12844
rect 7064 12832 7070 12844
rect 8021 12835 8079 12841
rect 8021 12832 8033 12835
rect 7064 12804 8033 12832
rect 7064 12792 7070 12804
rect 8021 12801 8033 12804
rect 8067 12832 8079 12835
rect 8110 12832 8116 12844
rect 8067 12804 8116 12832
rect 8067 12801 8079 12804
rect 8021 12795 8079 12801
rect 8110 12792 8116 12804
rect 8168 12792 8174 12844
rect 8288 12835 8346 12841
rect 8288 12801 8300 12835
rect 8334 12832 8346 12835
rect 8846 12832 8852 12844
rect 8334 12804 8852 12832
rect 8334 12801 8346 12804
rect 8288 12795 8346 12801
rect 8846 12792 8852 12804
rect 8904 12792 8910 12844
rect 9950 12832 9956 12844
rect 9911 12804 9956 12832
rect 9950 12792 9956 12804
rect 10008 12792 10014 12844
rect 10045 12835 10103 12841
rect 10045 12801 10057 12835
rect 10091 12801 10103 12835
rect 10045 12795 10103 12801
rect 10965 12835 11023 12841
rect 10965 12801 10977 12835
rect 11011 12832 11023 12835
rect 11606 12832 11612 12844
rect 11011 12804 11612 12832
rect 11011 12801 11023 12804
rect 10965 12795 11023 12801
rect 9674 12764 9680 12776
rect 9416 12736 9680 12764
rect 9416 12705 9444 12736
rect 9674 12724 9680 12736
rect 9732 12764 9738 12776
rect 10060 12764 10088 12795
rect 11606 12792 11612 12804
rect 11664 12792 11670 12844
rect 11784 12835 11842 12841
rect 11784 12801 11796 12835
rect 11830 12832 11842 12835
rect 12342 12832 12348 12844
rect 11830 12804 12348 12832
rect 11830 12801 11842 12804
rect 11784 12795 11842 12801
rect 12342 12792 12348 12804
rect 12400 12792 12406 12844
rect 14734 12792 14740 12844
rect 14792 12832 14798 12844
rect 15197 12835 15255 12841
rect 15197 12832 15209 12835
rect 14792 12804 15209 12832
rect 14792 12792 14798 12804
rect 15197 12801 15209 12804
rect 15243 12801 15255 12835
rect 15470 12832 15476 12844
rect 15431 12804 15476 12832
rect 15197 12795 15255 12801
rect 15470 12792 15476 12804
rect 15528 12792 15534 12844
rect 11514 12764 11520 12776
rect 9732 12736 10088 12764
rect 11475 12736 11520 12764
rect 9732 12724 9738 12736
rect 11514 12724 11520 12736
rect 11572 12724 11578 12776
rect 13170 12724 13176 12776
rect 13228 12764 13234 12776
rect 13357 12767 13415 12773
rect 13357 12764 13369 12767
rect 13228 12736 13369 12764
rect 13228 12724 13234 12736
rect 13357 12733 13369 12736
rect 13403 12733 13415 12767
rect 13357 12727 13415 12733
rect 14550 12724 14556 12776
rect 14608 12764 14614 12776
rect 15381 12767 15439 12773
rect 15381 12764 15393 12767
rect 14608 12736 15393 12764
rect 14608 12724 14614 12736
rect 15381 12733 15393 12736
rect 15427 12764 15439 12767
rect 15654 12764 15660 12776
rect 15427 12736 15660 12764
rect 15427 12733 15439 12736
rect 15381 12727 15439 12733
rect 15654 12724 15660 12736
rect 15712 12724 15718 12776
rect 9401 12699 9459 12705
rect 9401 12665 9413 12699
rect 9447 12665 9459 12699
rect 9401 12659 9459 12665
rect 10781 12699 10839 12705
rect 10781 12665 10793 12699
rect 10827 12696 10839 12699
rect 11054 12696 11060 12708
rect 10827 12668 11060 12696
rect 10827 12665 10839 12668
rect 10781 12659 10839 12665
rect 11054 12656 11060 12668
rect 11112 12656 11118 12708
rect 9674 12588 9680 12640
rect 9732 12628 9738 12640
rect 10229 12631 10287 12637
rect 10229 12628 10241 12631
rect 9732 12600 10241 12628
rect 9732 12588 9738 12600
rect 10229 12597 10241 12600
rect 10275 12597 10287 12631
rect 10229 12591 10287 12597
rect 12897 12631 12955 12637
rect 12897 12597 12909 12631
rect 12943 12628 12955 12631
rect 13262 12628 13268 12640
rect 12943 12600 13268 12628
rect 12943 12597 12955 12600
rect 12897 12591 12955 12597
rect 13262 12588 13268 12600
rect 13320 12628 13326 12640
rect 14550 12628 14556 12640
rect 13320 12600 14556 12628
rect 13320 12588 13326 12600
rect 14550 12588 14556 12600
rect 14608 12588 14614 12640
rect 14734 12628 14740 12640
rect 14695 12600 14740 12628
rect 14734 12588 14740 12600
rect 14792 12588 14798 12640
rect 15473 12631 15531 12637
rect 15473 12597 15485 12631
rect 15519 12628 15531 12631
rect 15562 12628 15568 12640
rect 15519 12600 15568 12628
rect 15519 12597 15531 12600
rect 15473 12591 15531 12597
rect 15562 12588 15568 12600
rect 15620 12588 15626 12640
rect 15755 12628 15783 12872
rect 17558 12869 17570 12872
rect 17604 12869 17616 12903
rect 17558 12863 17616 12869
rect 18138 12860 18144 12912
rect 18196 12900 18202 12912
rect 20898 12900 20904 12912
rect 18196 12872 20904 12900
rect 18196 12860 18202 12872
rect 20898 12860 20904 12872
rect 20956 12860 20962 12912
rect 26234 12900 26240 12912
rect 22066 12872 22416 12900
rect 16853 12835 16911 12841
rect 16853 12801 16865 12835
rect 16899 12832 16911 12835
rect 16942 12832 16948 12844
rect 16899 12804 16948 12832
rect 16899 12801 16911 12804
rect 16853 12795 16911 12801
rect 16942 12792 16948 12804
rect 17000 12792 17006 12844
rect 19981 12835 20039 12841
rect 19981 12801 19993 12835
rect 20027 12832 20039 12835
rect 20622 12832 20628 12844
rect 20027 12804 20628 12832
rect 20027 12801 20039 12804
rect 19981 12795 20039 12801
rect 20622 12792 20628 12804
rect 20680 12792 20686 12844
rect 16758 12724 16764 12776
rect 16816 12764 16822 12776
rect 17310 12764 17316 12776
rect 16816 12736 17316 12764
rect 16816 12724 16822 12736
rect 17310 12724 17316 12736
rect 17368 12724 17374 12776
rect 18598 12724 18604 12776
rect 18656 12764 18662 12776
rect 20165 12767 20223 12773
rect 20165 12764 20177 12767
rect 18656 12736 20177 12764
rect 18656 12724 18662 12736
rect 20165 12733 20177 12736
rect 20211 12764 20223 12767
rect 22066 12764 22094 12872
rect 22186 12832 22192 12844
rect 22147 12804 22192 12832
rect 22186 12792 22192 12804
rect 22244 12792 22250 12844
rect 22388 12773 22416 12872
rect 25976 12872 26240 12900
rect 23658 12832 23664 12844
rect 23619 12804 23664 12832
rect 23658 12792 23664 12804
rect 23716 12792 23722 12844
rect 24118 12832 24124 12844
rect 24079 12804 24124 12832
rect 24118 12792 24124 12804
rect 24176 12792 24182 12844
rect 24946 12832 24952 12844
rect 24907 12804 24952 12832
rect 24946 12792 24952 12804
rect 25004 12792 25010 12844
rect 25976 12841 26004 12872
rect 26234 12860 26240 12872
rect 26292 12900 26298 12912
rect 27614 12900 27620 12912
rect 26292 12872 27016 12900
rect 26292 12860 26298 12872
rect 26988 12844 27016 12872
rect 27448 12872 27620 12900
rect 25041 12835 25099 12841
rect 25041 12801 25053 12835
rect 25087 12832 25099 12835
rect 25961 12835 26019 12841
rect 25087 12804 25820 12832
rect 25087 12801 25099 12804
rect 25041 12795 25099 12801
rect 25792 12776 25820 12804
rect 25961 12801 25973 12835
rect 26007 12801 26019 12835
rect 25961 12795 26019 12801
rect 26053 12835 26111 12841
rect 26053 12801 26065 12835
rect 26099 12801 26111 12835
rect 26053 12795 26111 12801
rect 26145 12835 26203 12841
rect 26145 12801 26157 12835
rect 26191 12801 26203 12835
rect 26145 12795 26203 12801
rect 26329 12835 26387 12841
rect 26329 12801 26341 12835
rect 26375 12801 26387 12835
rect 26329 12795 26387 12801
rect 20211 12736 22094 12764
rect 22373 12767 22431 12773
rect 20211 12733 20223 12736
rect 20165 12727 20223 12733
rect 22373 12733 22385 12767
rect 22419 12733 22431 12767
rect 22373 12727 22431 12733
rect 24210 12724 24216 12776
rect 24268 12764 24274 12776
rect 24762 12764 24768 12776
rect 24268 12736 24768 12764
rect 24268 12724 24274 12736
rect 24762 12724 24768 12736
rect 24820 12764 24826 12776
rect 24857 12767 24915 12773
rect 24857 12764 24869 12767
rect 24820 12736 24869 12764
rect 24820 12724 24826 12736
rect 24857 12733 24869 12736
rect 24903 12733 24915 12767
rect 24857 12727 24915 12733
rect 25133 12767 25191 12773
rect 25133 12733 25145 12767
rect 25179 12733 25191 12767
rect 25133 12727 25191 12733
rect 23477 12699 23535 12705
rect 23477 12696 23489 12699
rect 18248 12668 23489 12696
rect 18248 12628 18276 12668
rect 23477 12665 23489 12668
rect 23523 12665 23535 12699
rect 23477 12659 23535 12665
rect 24578 12656 24584 12708
rect 24636 12696 24642 12708
rect 25148 12696 25176 12727
rect 25774 12724 25780 12776
rect 25832 12764 25838 12776
rect 26068 12764 26096 12795
rect 25832 12736 26096 12764
rect 26160 12764 26188 12795
rect 26344 12764 26372 12795
rect 26418 12792 26424 12844
rect 26476 12832 26482 12844
rect 26970 12832 26976 12844
rect 26476 12804 26521 12832
rect 26931 12804 26976 12832
rect 26476 12792 26482 12804
rect 26970 12792 26976 12804
rect 27028 12792 27034 12844
rect 27154 12832 27160 12844
rect 27115 12804 27160 12832
rect 27154 12792 27160 12804
rect 27212 12792 27218 12844
rect 26510 12764 26516 12776
rect 26160 12736 26280 12764
rect 26344 12736 26516 12764
rect 25832 12724 25838 12736
rect 26252 12708 26280 12736
rect 26510 12724 26516 12736
rect 26568 12724 26574 12776
rect 26786 12724 26792 12776
rect 26844 12764 26850 12776
rect 27249 12767 27307 12773
rect 27249 12764 27261 12767
rect 26844 12736 27261 12764
rect 26844 12724 26850 12736
rect 27249 12733 27261 12736
rect 27295 12733 27307 12767
rect 27249 12727 27307 12733
rect 27341 12767 27399 12773
rect 27341 12733 27353 12767
rect 27387 12764 27399 12767
rect 27448 12764 27476 12872
rect 27614 12860 27620 12872
rect 27672 12860 27678 12912
rect 27709 12903 27767 12909
rect 27709 12869 27721 12903
rect 27755 12900 27767 12903
rect 27755 12872 28396 12900
rect 27755 12869 27767 12872
rect 27709 12863 27767 12869
rect 27525 12835 27583 12841
rect 27525 12801 27537 12835
rect 27571 12801 27583 12835
rect 28166 12832 28172 12844
rect 28127 12804 28172 12832
rect 27525 12795 27583 12801
rect 27387 12736 27476 12764
rect 27387 12733 27399 12736
rect 27341 12727 27399 12733
rect 24636 12668 25176 12696
rect 24636 12656 24642 12668
rect 18690 12628 18696 12640
rect 15755 12600 18276 12628
rect 18651 12600 18696 12628
rect 18690 12588 18696 12600
rect 18748 12588 18754 12640
rect 19334 12588 19340 12640
rect 19392 12628 19398 12640
rect 19613 12631 19671 12637
rect 19613 12628 19625 12631
rect 19392 12600 19625 12628
rect 19392 12588 19398 12600
rect 19613 12597 19625 12600
rect 19659 12597 19671 12631
rect 21818 12628 21824 12640
rect 21779 12600 21824 12628
rect 19613 12591 19671 12597
rect 21818 12588 21824 12600
rect 21876 12588 21882 12640
rect 24673 12631 24731 12637
rect 24673 12597 24685 12631
rect 24719 12628 24731 12631
rect 24762 12628 24768 12640
rect 24719 12600 24768 12628
rect 24719 12597 24731 12600
rect 24673 12591 24731 12597
rect 24762 12588 24768 12600
rect 24820 12588 24826 12640
rect 25148 12628 25176 12668
rect 26234 12656 26240 12708
rect 26292 12696 26298 12708
rect 27540 12696 27568 12795
rect 28166 12792 28172 12804
rect 28224 12792 28230 12844
rect 28368 12841 28396 12872
rect 28353 12835 28411 12841
rect 28353 12801 28365 12835
rect 28399 12801 28411 12835
rect 37826 12832 37832 12844
rect 37787 12804 37832 12832
rect 28353 12795 28411 12801
rect 37826 12792 37832 12804
rect 37884 12792 37890 12844
rect 26292 12668 27568 12696
rect 28445 12699 28503 12705
rect 26292 12656 26298 12668
rect 28445 12665 28457 12699
rect 28491 12696 28503 12699
rect 38194 12696 38200 12708
rect 28491 12668 38200 12696
rect 28491 12665 28503 12668
rect 28445 12659 28503 12665
rect 38194 12656 38200 12668
rect 38252 12656 38258 12708
rect 26252 12628 26280 12656
rect 38010 12628 38016 12640
rect 25148 12600 26280 12628
rect 37971 12600 38016 12628
rect 38010 12588 38016 12600
rect 38068 12588 38074 12640
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 8846 12384 8852 12436
rect 8904 12424 8910 12436
rect 8941 12427 8999 12433
rect 8941 12424 8953 12427
rect 8904 12396 8953 12424
rect 8904 12384 8910 12396
rect 8941 12393 8953 12396
rect 8987 12393 8999 12427
rect 10962 12424 10968 12436
rect 10923 12396 10968 12424
rect 8941 12387 8999 12393
rect 10962 12384 10968 12396
rect 11020 12384 11026 12436
rect 12434 12384 12440 12436
rect 12492 12424 12498 12436
rect 13081 12427 13139 12433
rect 13081 12424 13093 12427
rect 12492 12396 13093 12424
rect 12492 12384 12498 12396
rect 13081 12393 13093 12396
rect 13127 12393 13139 12427
rect 13081 12387 13139 12393
rect 14734 12384 14740 12436
rect 14792 12424 14798 12436
rect 15105 12427 15163 12433
rect 15105 12424 15117 12427
rect 14792 12396 15117 12424
rect 14792 12384 14798 12396
rect 15105 12393 15117 12396
rect 15151 12393 15163 12427
rect 15286 12424 15292 12436
rect 15247 12396 15292 12424
rect 15105 12387 15163 12393
rect 15286 12384 15292 12396
rect 15344 12384 15350 12436
rect 17218 12424 17224 12436
rect 17179 12396 17224 12424
rect 17218 12384 17224 12396
rect 17276 12384 17282 12436
rect 17957 12427 18015 12433
rect 17957 12393 17969 12427
rect 18003 12424 18015 12427
rect 19426 12424 19432 12436
rect 18003 12396 19432 12424
rect 18003 12393 18015 12396
rect 17957 12387 18015 12393
rect 19426 12384 19432 12396
rect 19484 12384 19490 12436
rect 20622 12424 20628 12436
rect 20583 12396 20628 12424
rect 20622 12384 20628 12396
rect 20680 12384 20686 12436
rect 27433 12427 27491 12433
rect 27433 12393 27445 12427
rect 27479 12424 27491 12427
rect 27614 12424 27620 12436
rect 27479 12396 27620 12424
rect 27479 12393 27491 12396
rect 27433 12387 27491 12393
rect 27614 12384 27620 12396
rect 27672 12424 27678 12436
rect 28166 12424 28172 12436
rect 27672 12396 28172 12424
rect 27672 12384 27678 12396
rect 28166 12384 28172 12396
rect 28224 12384 28230 12436
rect 11606 12316 11612 12368
rect 11664 12356 11670 12368
rect 12621 12359 12679 12365
rect 12621 12356 12633 12359
rect 11664 12328 12633 12356
rect 11664 12316 11670 12328
rect 12621 12325 12633 12328
rect 12667 12325 12679 12359
rect 15194 12356 15200 12368
rect 12621 12319 12679 12325
rect 14016 12328 15200 12356
rect 8110 12248 8116 12300
rect 8168 12288 8174 12300
rect 9585 12291 9643 12297
rect 9585 12288 9597 12291
rect 8168 12260 9597 12288
rect 8168 12248 8174 12260
rect 9585 12257 9597 12260
rect 9631 12257 9643 12291
rect 9585 12251 9643 12257
rect 11425 12291 11483 12297
rect 11425 12257 11437 12291
rect 11471 12288 11483 12291
rect 11790 12288 11796 12300
rect 11471 12260 11796 12288
rect 11471 12257 11483 12260
rect 11425 12251 11483 12257
rect 11790 12248 11796 12260
rect 11848 12248 11854 12300
rect 12250 12288 12256 12300
rect 12211 12260 12256 12288
rect 12250 12248 12256 12260
rect 12308 12248 12314 12300
rect 14016 12288 14044 12328
rect 15194 12316 15200 12328
rect 15252 12356 15258 12368
rect 15252 12328 16068 12356
rect 15252 12316 15258 12328
rect 12452 12260 14044 12288
rect 14093 12291 14151 12297
rect 9122 12220 9128 12232
rect 9083 12192 9128 12220
rect 9122 12180 9128 12192
rect 9180 12180 9186 12232
rect 12452 12229 12480 12260
rect 14093 12257 14105 12291
rect 14139 12288 14151 12291
rect 14734 12288 14740 12300
rect 14139 12260 14740 12288
rect 14139 12257 14151 12260
rect 14093 12251 14151 12257
rect 14734 12248 14740 12260
rect 14792 12248 14798 12300
rect 16040 12297 16068 12328
rect 16025 12291 16083 12297
rect 16025 12257 16037 12291
rect 16071 12257 16083 12291
rect 18414 12288 18420 12300
rect 18375 12260 18420 12288
rect 16025 12251 16083 12257
rect 18414 12248 18420 12260
rect 18472 12248 18478 12300
rect 18598 12288 18604 12300
rect 18559 12260 18604 12288
rect 18598 12248 18604 12260
rect 18656 12248 18662 12300
rect 18690 12248 18696 12300
rect 18748 12288 18754 12300
rect 20640 12288 20668 12384
rect 25406 12356 25412 12368
rect 22388 12328 25412 12356
rect 22388 12297 22416 12328
rect 22373 12291 22431 12297
rect 18748 12260 19380 12288
rect 20640 12260 22140 12288
rect 18748 12248 18754 12260
rect 11609 12223 11667 12229
rect 11609 12189 11621 12223
rect 11655 12189 11667 12223
rect 11609 12183 11667 12189
rect 12437 12223 12495 12229
rect 12437 12189 12449 12223
rect 12483 12189 12495 12223
rect 12437 12183 12495 12189
rect 13265 12223 13323 12229
rect 13265 12189 13277 12223
rect 13311 12189 13323 12223
rect 13265 12183 13323 12189
rect 9490 12112 9496 12164
rect 9548 12152 9554 12164
rect 9830 12155 9888 12161
rect 9830 12152 9842 12155
rect 9548 12124 9842 12152
rect 9548 12112 9554 12124
rect 9830 12121 9842 12124
rect 9876 12121 9888 12155
rect 9830 12115 9888 12121
rect 11238 12112 11244 12164
rect 11296 12152 11302 12164
rect 11624 12152 11652 12183
rect 11296 12124 11652 12152
rect 11793 12155 11851 12161
rect 11296 12112 11302 12124
rect 11793 12121 11805 12155
rect 11839 12152 11851 12155
rect 13280 12152 13308 12183
rect 13446 12180 13452 12232
rect 13504 12220 13510 12232
rect 14277 12223 14335 12229
rect 14277 12220 14289 12223
rect 13504 12192 14289 12220
rect 13504 12180 13510 12192
rect 14277 12189 14289 12192
rect 14323 12189 14335 12223
rect 14277 12183 14335 12189
rect 14642 12180 14648 12232
rect 14700 12220 14706 12232
rect 15749 12223 15807 12229
rect 15749 12220 15761 12223
rect 14700 12192 15761 12220
rect 14700 12180 14706 12192
rect 15749 12189 15761 12192
rect 15795 12189 15807 12223
rect 15749 12183 15807 12189
rect 18325 12223 18383 12229
rect 18325 12189 18337 12223
rect 18371 12220 18383 12223
rect 18708 12220 18736 12248
rect 18371 12192 18736 12220
rect 19245 12223 19303 12229
rect 18371 12189 18383 12192
rect 18325 12183 18383 12189
rect 19245 12189 19257 12223
rect 19291 12189 19303 12223
rect 19352 12220 19380 12260
rect 21269 12223 21327 12229
rect 19352 12192 21220 12220
rect 19245 12183 19303 12189
rect 11839 12124 13308 12152
rect 11839 12121 11851 12124
rect 11793 12115 11851 12121
rect 14550 12112 14556 12164
rect 14608 12152 14614 12164
rect 14921 12155 14979 12161
rect 14921 12152 14933 12155
rect 14608 12124 14933 12152
rect 14608 12112 14614 12124
rect 14921 12121 14933 12124
rect 14967 12152 14979 12155
rect 15470 12152 15476 12164
rect 14967 12124 15476 12152
rect 14967 12121 14979 12124
rect 14921 12115 14979 12121
rect 15470 12112 15476 12124
rect 15528 12112 15534 12164
rect 15764 12152 15792 12183
rect 16482 12152 16488 12164
rect 15764 12124 16488 12152
rect 16482 12112 16488 12124
rect 16540 12152 16546 12164
rect 17129 12155 17187 12161
rect 17129 12152 17141 12155
rect 16540 12124 17141 12152
rect 16540 12112 16546 12124
rect 17129 12121 17141 12124
rect 17175 12121 17187 12155
rect 17129 12115 17187 12121
rect 17310 12112 17316 12164
rect 17368 12152 17374 12164
rect 19260 12152 19288 12183
rect 19512 12155 19570 12161
rect 17368 12124 19334 12152
rect 17368 12112 17374 12124
rect 14274 12044 14280 12096
rect 14332 12084 14338 12096
rect 14461 12087 14519 12093
rect 14461 12084 14473 12087
rect 14332 12056 14473 12084
rect 14332 12044 14338 12056
rect 14461 12053 14473 12056
rect 14507 12053 14519 12087
rect 14461 12047 14519 12053
rect 14734 12044 14740 12096
rect 14792 12084 14798 12096
rect 15121 12087 15179 12093
rect 15121 12084 15133 12087
rect 14792 12056 15133 12084
rect 14792 12044 14798 12056
rect 15121 12053 15133 12056
rect 15167 12053 15179 12087
rect 19306 12084 19334 12124
rect 19512 12121 19524 12155
rect 19558 12152 19570 12155
rect 21192 12152 21220 12192
rect 21269 12189 21281 12223
rect 21315 12220 21327 12223
rect 21358 12220 21364 12232
rect 21315 12192 21364 12220
rect 21315 12189 21327 12192
rect 21269 12183 21327 12189
rect 21358 12180 21364 12192
rect 21416 12180 21422 12232
rect 22112 12229 22140 12260
rect 22373 12257 22385 12291
rect 22419 12257 22431 12291
rect 23382 12288 23388 12300
rect 23343 12260 23388 12288
rect 22373 12251 22431 12257
rect 23382 12248 23388 12260
rect 23440 12248 23446 12300
rect 23492 12297 23520 12328
rect 25406 12316 25412 12328
rect 25464 12316 25470 12368
rect 26234 12316 26240 12368
rect 26292 12316 26298 12368
rect 23477 12291 23535 12297
rect 23477 12257 23489 12291
rect 23523 12257 23535 12291
rect 23477 12251 23535 12257
rect 23750 12248 23756 12300
rect 23808 12288 23814 12300
rect 24578 12288 24584 12300
rect 23808 12260 24584 12288
rect 23808 12248 23814 12260
rect 24578 12248 24584 12260
rect 24636 12288 24642 12300
rect 24673 12291 24731 12297
rect 24673 12288 24685 12291
rect 24636 12260 24685 12288
rect 24636 12248 24642 12260
rect 24673 12257 24685 12260
rect 24719 12257 24731 12291
rect 26252 12288 26280 12316
rect 26252 12260 26372 12288
rect 24673 12251 24731 12257
rect 22097 12223 22155 12229
rect 22097 12189 22109 12223
rect 22143 12189 22155 12223
rect 22097 12183 22155 12189
rect 22186 12180 22192 12232
rect 22244 12220 22250 12232
rect 23293 12223 23351 12229
rect 23293 12220 23305 12223
rect 22244 12192 23305 12220
rect 22244 12180 22250 12192
rect 23293 12189 23305 12192
rect 23339 12189 23351 12223
rect 23293 12183 23351 12189
rect 23566 12180 23572 12232
rect 23624 12220 23630 12232
rect 24397 12223 24455 12229
rect 24397 12220 24409 12223
rect 23624 12192 24409 12220
rect 23624 12180 23630 12192
rect 24397 12189 24409 12192
rect 24443 12189 24455 12223
rect 24397 12183 24455 12189
rect 25866 12180 25872 12232
rect 25924 12220 25930 12232
rect 26344 12229 26372 12260
rect 26620 12260 27292 12288
rect 26620 12232 26648 12260
rect 26237 12223 26295 12229
rect 26237 12220 26249 12223
rect 25924 12192 26249 12220
rect 25924 12180 25930 12192
rect 26237 12189 26249 12192
rect 26283 12189 26295 12223
rect 26237 12183 26295 12189
rect 26329 12223 26387 12229
rect 26329 12189 26341 12223
rect 26375 12189 26387 12223
rect 26329 12183 26387 12189
rect 26418 12180 26424 12232
rect 26476 12220 26482 12232
rect 26513 12223 26571 12229
rect 26513 12220 26525 12223
rect 26476 12192 26525 12220
rect 26476 12180 26482 12192
rect 26513 12189 26525 12192
rect 26559 12189 26571 12223
rect 26513 12183 26571 12189
rect 26602 12180 26608 12232
rect 26660 12220 26666 12232
rect 27062 12220 27068 12232
rect 26660 12192 26705 12220
rect 27023 12192 27068 12220
rect 26660 12180 26666 12192
rect 27062 12180 27068 12192
rect 27120 12180 27126 12232
rect 27264 12229 27292 12260
rect 27249 12223 27307 12229
rect 27249 12189 27261 12223
rect 27295 12189 27307 12223
rect 27249 12183 27307 12189
rect 26053 12155 26111 12161
rect 19558 12124 21128 12152
rect 21192 12124 22232 12152
rect 19558 12121 19570 12124
rect 19512 12115 19570 12121
rect 20714 12084 20720 12096
rect 19306 12056 20720 12084
rect 15121 12047 15179 12053
rect 20714 12044 20720 12056
rect 20772 12084 20778 12096
rect 20990 12084 20996 12096
rect 20772 12056 20996 12084
rect 20772 12044 20778 12056
rect 20990 12044 20996 12056
rect 21048 12044 21054 12096
rect 21100 12093 21128 12124
rect 21085 12087 21143 12093
rect 21085 12053 21097 12087
rect 21131 12053 21143 12087
rect 21726 12084 21732 12096
rect 21687 12056 21732 12084
rect 21085 12047 21143 12053
rect 21726 12044 21732 12056
rect 21784 12044 21790 12096
rect 22204 12093 22232 12124
rect 26053 12121 26065 12155
rect 26099 12152 26111 12155
rect 37826 12152 37832 12164
rect 26099 12124 37832 12152
rect 26099 12121 26111 12124
rect 26053 12115 26111 12121
rect 37826 12112 37832 12124
rect 37884 12112 37890 12164
rect 22189 12087 22247 12093
rect 22189 12053 22201 12087
rect 22235 12053 22247 12087
rect 22189 12047 22247 12053
rect 22738 12044 22744 12096
rect 22796 12084 22802 12096
rect 22925 12087 22983 12093
rect 22925 12084 22937 12087
rect 22796 12056 22937 12084
rect 22796 12044 22802 12056
rect 22925 12053 22937 12056
rect 22971 12053 22983 12087
rect 22925 12047 22983 12053
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 9490 11880 9496 11892
rect 9451 11852 9496 11880
rect 9490 11840 9496 11852
rect 9548 11840 9554 11892
rect 14093 11883 14151 11889
rect 14093 11849 14105 11883
rect 14139 11849 14151 11883
rect 14093 11843 14151 11849
rect 19521 11883 19579 11889
rect 19521 11849 19533 11883
rect 19567 11880 19579 11883
rect 21358 11880 21364 11892
rect 19567 11852 21364 11880
rect 19567 11849 19579 11852
rect 19521 11843 19579 11849
rect 14108 11812 14136 11843
rect 21358 11840 21364 11852
rect 21416 11840 21422 11892
rect 27065 11883 27123 11889
rect 27065 11849 27077 11883
rect 27111 11880 27123 11883
rect 27154 11880 27160 11892
rect 27111 11852 27160 11880
rect 27111 11849 27123 11852
rect 27065 11843 27123 11849
rect 27154 11840 27160 11852
rect 27212 11840 27218 11892
rect 14982 11815 15040 11821
rect 14982 11812 14994 11815
rect 14108 11784 14994 11812
rect 14982 11781 14994 11784
rect 15028 11781 15040 11815
rect 21818 11812 21824 11824
rect 14982 11775 15040 11781
rect 20180 11784 21824 11812
rect 8662 11744 8668 11756
rect 8623 11716 8668 11744
rect 8662 11704 8668 11716
rect 8720 11704 8726 11756
rect 9674 11744 9680 11756
rect 9635 11716 9680 11744
rect 9674 11704 9680 11716
rect 9732 11704 9738 11756
rect 10137 11747 10195 11753
rect 10137 11713 10149 11747
rect 10183 11744 10195 11747
rect 11517 11747 11575 11753
rect 10183 11716 11468 11744
rect 10183 11713 10195 11716
rect 10137 11707 10195 11713
rect 8202 11636 8208 11688
rect 8260 11676 8266 11688
rect 10318 11676 10324 11688
rect 8260 11648 10324 11676
rect 8260 11636 8266 11648
rect 10318 11636 10324 11648
rect 10376 11676 10382 11688
rect 10413 11679 10471 11685
rect 10413 11676 10425 11679
rect 10376 11648 10425 11676
rect 10376 11636 10382 11648
rect 10413 11645 10425 11648
rect 10459 11645 10471 11679
rect 11440 11676 11468 11716
rect 11517 11713 11529 11747
rect 11563 11744 11575 11747
rect 12618 11744 12624 11756
rect 11563 11716 12624 11744
rect 11563 11713 11575 11716
rect 11517 11707 11575 11713
rect 12618 11704 12624 11716
rect 12676 11744 12682 11756
rect 12894 11744 12900 11756
rect 12676 11716 12900 11744
rect 12676 11704 12682 11716
rect 12894 11704 12900 11716
rect 12952 11704 12958 11756
rect 13081 11747 13139 11753
rect 13081 11713 13093 11747
rect 13127 11744 13139 11747
rect 13446 11744 13452 11756
rect 13127 11716 13452 11744
rect 13127 11713 13139 11716
rect 13081 11707 13139 11713
rect 13446 11704 13452 11716
rect 13504 11704 13510 11756
rect 14274 11744 14280 11756
rect 14235 11716 14280 11744
rect 14274 11704 14280 11716
rect 14332 11704 14338 11756
rect 14737 11747 14795 11753
rect 14737 11713 14749 11747
rect 14783 11744 14795 11747
rect 14826 11744 14832 11756
rect 14783 11716 14832 11744
rect 14783 11713 14795 11716
rect 14737 11707 14795 11713
rect 14826 11704 14832 11716
rect 14884 11704 14890 11756
rect 16482 11704 16488 11756
rect 16540 11744 16546 11756
rect 16945 11747 17003 11753
rect 16945 11744 16957 11747
rect 16540 11716 16957 11744
rect 16540 11704 16546 11716
rect 16945 11713 16957 11716
rect 16991 11744 17003 11747
rect 18049 11747 18107 11753
rect 18049 11744 18061 11747
rect 16991 11716 18061 11744
rect 16991 11713 17003 11716
rect 16945 11707 17003 11713
rect 18049 11713 18061 11716
rect 18095 11713 18107 11747
rect 19334 11744 19340 11756
rect 19295 11716 19340 11744
rect 18049 11707 18107 11713
rect 19334 11704 19340 11716
rect 19392 11704 19398 11756
rect 20180 11753 20208 11784
rect 21818 11772 21824 11784
rect 21876 11772 21882 11824
rect 20165 11747 20223 11753
rect 20165 11713 20177 11747
rect 20211 11713 20223 11747
rect 20165 11707 20223 11713
rect 20349 11747 20407 11753
rect 20349 11713 20361 11747
rect 20395 11744 20407 11747
rect 20993 11747 21051 11753
rect 20993 11744 21005 11747
rect 20395 11716 21005 11744
rect 20395 11713 20407 11716
rect 20349 11707 20407 11713
rect 20993 11713 21005 11716
rect 21039 11713 21051 11747
rect 20993 11707 21051 11713
rect 21726 11704 21732 11756
rect 21784 11744 21790 11756
rect 22925 11747 22983 11753
rect 22925 11744 22937 11747
rect 21784 11716 22937 11744
rect 21784 11704 21790 11716
rect 22925 11713 22937 11716
rect 22971 11744 22983 11747
rect 23474 11744 23480 11756
rect 22971 11716 23480 11744
rect 22971 11713 22983 11716
rect 22925 11707 22983 11713
rect 23474 11704 23480 11716
rect 23532 11744 23538 11756
rect 23661 11747 23719 11753
rect 23661 11744 23673 11747
rect 23532 11716 23673 11744
rect 23532 11704 23538 11716
rect 23661 11713 23673 11716
rect 23707 11713 23719 11747
rect 24949 11747 25007 11753
rect 24949 11744 24961 11747
rect 23661 11707 23719 11713
rect 23860 11716 24961 11744
rect 12805 11679 12863 11685
rect 12805 11676 12817 11679
rect 11440 11648 12817 11676
rect 10413 11639 10471 11645
rect 12805 11645 12817 11648
rect 12851 11676 12863 11679
rect 14642 11676 14648 11688
rect 12851 11648 14648 11676
rect 12851 11645 12863 11648
rect 12805 11639 12863 11645
rect 14642 11636 14648 11648
rect 14700 11636 14706 11688
rect 16114 11636 16120 11688
rect 16172 11676 16178 11688
rect 16669 11679 16727 11685
rect 16669 11676 16681 11679
rect 16172 11648 16681 11676
rect 16172 11636 16178 11648
rect 16669 11645 16681 11648
rect 16715 11645 16727 11679
rect 16669 11639 16727 11645
rect 19153 11679 19211 11685
rect 19153 11645 19165 11679
rect 19199 11676 19211 11679
rect 19242 11676 19248 11688
rect 19199 11648 19248 11676
rect 19199 11645 19211 11648
rect 19153 11639 19211 11645
rect 19242 11636 19248 11648
rect 19300 11676 19306 11688
rect 19981 11679 20039 11685
rect 19981 11676 19993 11679
rect 19300 11648 19993 11676
rect 19300 11636 19306 11648
rect 19981 11645 19993 11648
rect 20027 11645 20039 11679
rect 22738 11676 22744 11688
rect 22699 11648 22744 11676
rect 19981 11639 20039 11645
rect 22738 11636 22744 11648
rect 22796 11676 22802 11688
rect 23566 11676 23572 11688
rect 22796 11648 23572 11676
rect 22796 11636 22802 11648
rect 23566 11636 23572 11648
rect 23624 11676 23630 11688
rect 23860 11676 23888 11716
rect 24949 11713 24961 11716
rect 24995 11713 25007 11747
rect 25869 11747 25927 11753
rect 25869 11744 25881 11747
rect 24949 11707 25007 11713
rect 25424 11716 25881 11744
rect 23624 11648 23888 11676
rect 23937 11679 23995 11685
rect 23624 11636 23630 11648
rect 23937 11645 23949 11679
rect 23983 11676 23995 11679
rect 24210 11676 24216 11688
rect 23983 11648 24216 11676
rect 23983 11645 23995 11648
rect 23937 11639 23995 11645
rect 24210 11636 24216 11648
rect 24268 11636 24274 11688
rect 25424 11685 25452 11716
rect 25869 11713 25881 11716
rect 25915 11744 25927 11747
rect 26050 11744 26056 11756
rect 25915 11716 26056 11744
rect 25915 11713 25927 11716
rect 25869 11707 25927 11713
rect 26050 11704 26056 11716
rect 26108 11704 26114 11756
rect 26418 11704 26424 11756
rect 26476 11744 26482 11756
rect 26973 11747 27031 11753
rect 26973 11744 26985 11747
rect 26476 11716 26985 11744
rect 26476 11704 26482 11716
rect 26973 11713 26985 11716
rect 27019 11744 27031 11747
rect 27062 11744 27068 11756
rect 27019 11716 27068 11744
rect 27019 11713 27031 11716
rect 26973 11707 27031 11713
rect 27062 11704 27068 11716
rect 27120 11704 27126 11756
rect 27614 11744 27620 11756
rect 27575 11716 27620 11744
rect 27614 11704 27620 11716
rect 27672 11704 27678 11756
rect 25409 11679 25467 11685
rect 25409 11645 25421 11679
rect 25455 11645 25467 11679
rect 25958 11676 25964 11688
rect 25919 11648 25964 11676
rect 25409 11639 25467 11645
rect 25958 11636 25964 11648
rect 26016 11636 26022 11688
rect 26234 11636 26240 11688
rect 26292 11676 26298 11688
rect 27709 11679 27767 11685
rect 27709 11676 27721 11679
rect 26292 11648 27721 11676
rect 26292 11636 26298 11648
rect 27709 11645 27721 11648
rect 27755 11645 27767 11679
rect 27709 11639 27767 11645
rect 18233 11611 18291 11617
rect 18233 11577 18245 11611
rect 18279 11608 18291 11611
rect 21910 11608 21916 11620
rect 18279 11580 21916 11608
rect 18279 11577 18291 11580
rect 18233 11571 18291 11577
rect 21910 11568 21916 11580
rect 21968 11568 21974 11620
rect 26786 11608 26792 11620
rect 24136 11580 26792 11608
rect 24136 11552 24164 11580
rect 26786 11568 26792 11580
rect 26844 11568 26850 11620
rect 8481 11543 8539 11549
rect 8481 11509 8493 11543
rect 8527 11540 8539 11543
rect 9030 11540 9036 11552
rect 8527 11512 9036 11540
rect 8527 11509 8539 11512
rect 8481 11503 8539 11509
rect 9030 11500 9036 11512
rect 9088 11500 9094 11552
rect 11330 11500 11336 11552
rect 11388 11540 11394 11552
rect 11701 11543 11759 11549
rect 11701 11540 11713 11543
rect 11388 11512 11713 11540
rect 11388 11500 11394 11512
rect 11701 11509 11713 11512
rect 11747 11540 11759 11543
rect 12158 11540 12164 11552
rect 11747 11512 12164 11540
rect 11747 11509 11759 11512
rect 11701 11503 11759 11509
rect 12158 11500 12164 11512
rect 12216 11500 12222 11552
rect 15470 11500 15476 11552
rect 15528 11540 15534 11552
rect 16117 11543 16175 11549
rect 16117 11540 16129 11543
rect 15528 11512 16129 11540
rect 15528 11500 15534 11512
rect 16117 11509 16129 11512
rect 16163 11509 16175 11543
rect 20806 11540 20812 11552
rect 20767 11512 20812 11540
rect 16117 11503 16175 11509
rect 20806 11500 20812 11512
rect 20864 11500 20870 11552
rect 23109 11543 23167 11549
rect 23109 11509 23121 11543
rect 23155 11540 23167 11543
rect 24118 11540 24124 11552
rect 23155 11512 24124 11540
rect 23155 11509 23167 11512
rect 23109 11503 23167 11509
rect 24118 11500 24124 11512
rect 24176 11500 24182 11552
rect 24210 11500 24216 11552
rect 24268 11540 24274 11552
rect 25041 11543 25099 11549
rect 25041 11540 25053 11543
rect 24268 11512 25053 11540
rect 24268 11500 24274 11512
rect 25041 11509 25053 11512
rect 25087 11509 25099 11543
rect 25041 11503 25099 11509
rect 25314 11500 25320 11552
rect 25372 11540 25378 11552
rect 25869 11543 25927 11549
rect 25869 11540 25881 11543
rect 25372 11512 25881 11540
rect 25372 11500 25378 11512
rect 25869 11509 25881 11512
rect 25915 11540 25927 11543
rect 26142 11540 26148 11552
rect 25915 11512 26148 11540
rect 25915 11509 25927 11512
rect 25869 11503 25927 11509
rect 26142 11500 26148 11512
rect 26200 11500 26206 11552
rect 26237 11543 26295 11549
rect 26237 11509 26249 11543
rect 26283 11540 26295 11543
rect 26326 11540 26332 11552
rect 26283 11512 26332 11540
rect 26283 11509 26295 11512
rect 26237 11503 26295 11509
rect 26326 11500 26332 11512
rect 26384 11500 26390 11552
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 12161 11339 12219 11345
rect 6886 11308 11744 11336
rect 1397 11135 1455 11141
rect 1397 11101 1409 11135
rect 1443 11132 1455 11135
rect 6886 11132 6914 11308
rect 11716 11268 11744 11308
rect 12161 11305 12173 11339
rect 12207 11336 12219 11339
rect 12250 11336 12256 11348
rect 12207 11308 12256 11336
rect 12207 11305 12219 11308
rect 12161 11299 12219 11305
rect 12250 11296 12256 11308
rect 12308 11296 12314 11348
rect 14734 11336 14740 11348
rect 12360 11308 14504 11336
rect 14695 11308 14740 11336
rect 12360 11268 12388 11308
rect 11716 11240 12388 11268
rect 14476 11268 14504 11308
rect 14734 11296 14740 11308
rect 14792 11296 14798 11348
rect 24949 11339 25007 11345
rect 24949 11336 24961 11339
rect 14844 11308 24961 11336
rect 14844 11268 14872 11308
rect 24949 11305 24961 11308
rect 24995 11305 25007 11339
rect 24949 11299 25007 11305
rect 14476 11240 14872 11268
rect 16301 11271 16359 11277
rect 16301 11237 16313 11271
rect 16347 11268 16359 11271
rect 18138 11268 18144 11280
rect 16347 11240 16804 11268
rect 18099 11240 18144 11268
rect 16347 11237 16359 11240
rect 16301 11231 16359 11237
rect 12894 11160 12900 11212
rect 12952 11200 12958 11212
rect 15473 11203 15531 11209
rect 15473 11200 15485 11203
rect 12952 11172 15485 11200
rect 12952 11160 12958 11172
rect 15473 11169 15485 11172
rect 15519 11169 15531 11203
rect 15473 11163 15531 11169
rect 15933 11203 15991 11209
rect 15933 11169 15945 11203
rect 15979 11200 15991 11203
rect 16666 11200 16672 11212
rect 15979 11172 16672 11200
rect 15979 11169 15991 11172
rect 15933 11163 15991 11169
rect 16666 11160 16672 11172
rect 16724 11160 16730 11212
rect 16776 11200 16804 11240
rect 18138 11228 18144 11240
rect 18196 11268 18202 11280
rect 18506 11268 18512 11280
rect 18196 11240 18512 11268
rect 18196 11228 18202 11240
rect 18506 11228 18512 11240
rect 18564 11228 18570 11280
rect 19245 11271 19303 11277
rect 19245 11237 19257 11271
rect 19291 11268 19303 11271
rect 19334 11268 19340 11280
rect 19291 11240 19340 11268
rect 19291 11237 19303 11240
rect 19245 11231 19303 11237
rect 19334 11228 19340 11240
rect 19392 11228 19398 11280
rect 22097 11271 22155 11277
rect 22097 11237 22109 11271
rect 22143 11268 22155 11271
rect 22186 11268 22192 11280
rect 22143 11240 22192 11268
rect 22143 11237 22155 11240
rect 22097 11231 22155 11237
rect 22186 11228 22192 11240
rect 22244 11228 22250 11280
rect 23845 11271 23903 11277
rect 23845 11237 23857 11271
rect 23891 11268 23903 11271
rect 24670 11268 24676 11280
rect 23891 11240 24676 11268
rect 23891 11237 23903 11240
rect 23845 11231 23903 11237
rect 24670 11228 24676 11240
rect 24728 11268 24734 11280
rect 26418 11268 26424 11280
rect 24728 11240 26424 11268
rect 24728 11228 24734 11240
rect 26418 11228 26424 11240
rect 26476 11228 26482 11280
rect 26789 11271 26847 11277
rect 26789 11237 26801 11271
rect 26835 11237 26847 11271
rect 26789 11231 26847 11237
rect 20714 11200 20720 11212
rect 16776 11172 16896 11200
rect 20675 11172 20720 11200
rect 1443 11104 6914 11132
rect 7009 11135 7067 11141
rect 1443 11101 1455 11104
rect 1397 11095 1455 11101
rect 7009 11101 7021 11135
rect 7055 11132 7067 11135
rect 8110 11132 8116 11144
rect 7055 11104 8116 11132
rect 7055 11101 7067 11104
rect 7009 11095 7067 11101
rect 8110 11092 8116 11104
rect 8168 11132 8174 11144
rect 8941 11135 8999 11141
rect 8941 11132 8953 11135
rect 8168 11104 8953 11132
rect 8168 11092 8174 11104
rect 8941 11101 8953 11104
rect 8987 11101 8999 11135
rect 8941 11095 8999 11101
rect 7276 11067 7334 11073
rect 7276 11033 7288 11067
rect 7322 11064 7334 11067
rect 7558 11064 7564 11076
rect 7322 11036 7564 11064
rect 7322 11033 7334 11036
rect 7276 11027 7334 11033
rect 7558 11024 7564 11036
rect 7616 11024 7622 11076
rect 8956 11064 8984 11095
rect 9030 11092 9036 11144
rect 9088 11132 9094 11144
rect 9197 11135 9255 11141
rect 9197 11132 9209 11135
rect 9088 11104 9209 11132
rect 9088 11092 9094 11104
rect 9197 11101 9209 11104
rect 9243 11101 9255 11135
rect 9197 11095 9255 11101
rect 10226 11092 10232 11144
rect 10284 11132 10290 11144
rect 10781 11135 10839 11141
rect 10781 11132 10793 11135
rect 10284 11104 10793 11132
rect 10284 11092 10290 11104
rect 10781 11101 10793 11104
rect 10827 11132 10839 11135
rect 10870 11132 10876 11144
rect 10827 11104 10876 11132
rect 10827 11101 10839 11104
rect 10781 11095 10839 11101
rect 10870 11092 10876 11104
rect 10928 11092 10934 11144
rect 13265 11135 13323 11141
rect 13265 11101 13277 11135
rect 13311 11101 13323 11135
rect 13265 11095 13323 11101
rect 13357 11135 13415 11141
rect 13357 11101 13369 11135
rect 13403 11132 13415 11135
rect 13446 11132 13452 11144
rect 13403 11104 13452 11132
rect 13403 11101 13415 11104
rect 13357 11095 13415 11101
rect 8956 11036 9260 11064
rect 1578 10996 1584 11008
rect 1539 10968 1584 10996
rect 1578 10956 1584 10968
rect 1636 10956 1642 11008
rect 8386 10996 8392 11008
rect 8347 10968 8392 10996
rect 8386 10956 8392 10968
rect 8444 10956 8450 11008
rect 9232 10996 9260 11036
rect 9306 11024 9312 11076
rect 9364 11064 9370 11076
rect 11054 11073 11060 11076
rect 9364 11036 10364 11064
rect 9364 11024 9370 11036
rect 10226 10996 10232 11008
rect 9232 10968 10232 10996
rect 10226 10956 10232 10968
rect 10284 10956 10290 11008
rect 10336 11005 10364 11036
rect 11048 11027 11060 11073
rect 11112 11064 11118 11076
rect 13280 11064 13308 11095
rect 13446 11092 13452 11104
rect 13504 11092 13510 11144
rect 13541 11135 13599 11141
rect 13541 11101 13553 11135
rect 13587 11132 13599 11135
rect 14274 11132 14280 11144
rect 13587 11104 14280 11132
rect 13587 11101 13599 11104
rect 13541 11095 13599 11101
rect 14274 11092 14280 11104
rect 14332 11092 14338 11144
rect 14366 11092 14372 11144
rect 14424 11132 14430 11144
rect 15289 11135 15347 11141
rect 14424 11104 14469 11132
rect 14424 11092 14430 11104
rect 15289 11101 15301 11135
rect 15335 11132 15347 11135
rect 16114 11132 16120 11144
rect 15335 11104 16120 11132
rect 15335 11101 15347 11104
rect 15289 11095 15347 11101
rect 16114 11092 16120 11104
rect 16172 11092 16178 11144
rect 16574 11092 16580 11144
rect 16632 11132 16638 11144
rect 16758 11132 16764 11144
rect 16632 11104 16764 11132
rect 16632 11092 16638 11104
rect 16758 11092 16764 11104
rect 16816 11092 16822 11144
rect 16868 11132 16896 11172
rect 20714 11160 20720 11172
rect 20772 11160 20778 11212
rect 25682 11200 25688 11212
rect 24412 11172 25688 11200
rect 18598 11132 18604 11144
rect 16868 11104 18604 11132
rect 18598 11092 18604 11104
rect 18656 11092 18662 11144
rect 19426 11132 19432 11144
rect 19387 11104 19432 11132
rect 19426 11092 19432 11104
rect 19484 11092 19490 11144
rect 20806 11092 20812 11144
rect 20864 11132 20870 11144
rect 20973 11135 21031 11141
rect 20973 11132 20985 11135
rect 20864 11104 20985 11132
rect 20864 11092 20870 11104
rect 20973 11101 20985 11104
rect 21019 11101 21031 11135
rect 23474 11132 23480 11144
rect 23435 11104 23480 11132
rect 20973 11095 21031 11101
rect 23474 11092 23480 11104
rect 23532 11092 23538 11144
rect 23566 11092 23572 11144
rect 23624 11132 23630 11144
rect 24412 11141 24440 11172
rect 25682 11160 25688 11172
rect 25740 11160 25746 11212
rect 26234 11200 26240 11212
rect 25792 11172 26240 11200
rect 23661 11135 23719 11141
rect 23661 11132 23673 11135
rect 23624 11104 23673 11132
rect 23624 11092 23630 11104
rect 23661 11101 23673 11104
rect 23707 11101 23719 11135
rect 23661 11095 23719 11101
rect 24397 11135 24455 11141
rect 24397 11101 24409 11135
rect 24443 11101 24455 11135
rect 24397 11095 24455 11101
rect 24762 11092 24768 11144
rect 24820 11141 24826 11144
rect 25792 11141 25820 11172
rect 26234 11160 26240 11172
rect 26292 11160 26298 11212
rect 26510 11200 26516 11212
rect 26344 11172 26516 11200
rect 26344 11141 26372 11172
rect 26510 11160 26516 11172
rect 26568 11160 26574 11212
rect 26602 11160 26608 11212
rect 26660 11200 26666 11212
rect 26804 11200 26832 11231
rect 26660 11172 26832 11200
rect 26660 11160 26666 11172
rect 24820 11132 24828 11141
rect 25777 11135 25835 11141
rect 24820 11104 24865 11132
rect 24820 11095 24828 11104
rect 25777 11101 25789 11135
rect 25823 11101 25835 11135
rect 25777 11095 25835 11101
rect 26329 11135 26387 11141
rect 26329 11101 26341 11135
rect 26375 11101 26387 11135
rect 26329 11095 26387 11101
rect 26421 11135 26479 11141
rect 26421 11101 26433 11135
rect 26467 11101 26479 11135
rect 26421 11095 26479 11101
rect 26697 11135 26755 11141
rect 26697 11101 26709 11135
rect 26743 11101 26755 11135
rect 26697 11095 26755 11101
rect 24820 11092 24826 11095
rect 14185 11067 14243 11073
rect 14185 11064 14197 11067
rect 11112 11036 11148 11064
rect 13280 11036 14197 11064
rect 11054 11024 11060 11027
rect 11112 11024 11118 11036
rect 14185 11033 14197 11036
rect 14231 11064 14243 11067
rect 15470 11064 15476 11076
rect 14231 11036 15476 11064
rect 14231 11033 14243 11036
rect 14185 11027 14243 11033
rect 15470 11024 15476 11036
rect 15528 11024 15534 11076
rect 16850 11024 16856 11076
rect 16908 11064 16914 11076
rect 17006 11067 17064 11073
rect 17006 11064 17018 11067
rect 16908 11036 17018 11064
rect 16908 11024 16914 11036
rect 17006 11033 17018 11036
rect 17052 11033 17064 11067
rect 24578 11064 24584 11076
rect 24539 11036 24584 11064
rect 17006 11027 17064 11033
rect 24578 11024 24584 11036
rect 24636 11024 24642 11076
rect 24673 11067 24731 11073
rect 24673 11033 24685 11067
rect 24719 11064 24731 11067
rect 25406 11064 25412 11076
rect 24719 11036 25412 11064
rect 24719 11033 24731 11036
rect 24673 11027 24731 11033
rect 25406 11024 25412 11036
rect 25464 11024 25470 11076
rect 25958 11024 25964 11076
rect 26016 11064 26022 11076
rect 26436 11064 26464 11095
rect 26712 11064 26740 11095
rect 26786 11092 26792 11144
rect 26844 11132 26850 11144
rect 26844 11104 26889 11132
rect 26844 11092 26850 11104
rect 26016 11036 26464 11064
rect 26528 11036 26740 11064
rect 26016 11024 26022 11036
rect 10321 10999 10379 11005
rect 10321 10965 10333 10999
rect 10367 10965 10379 10999
rect 10321 10959 10379 10965
rect 14090 10956 14096 11008
rect 14148 10996 14154 11008
rect 14461 10999 14519 11005
rect 14461 10996 14473 10999
rect 14148 10968 14473 10996
rect 14148 10956 14154 10968
rect 14461 10965 14473 10968
rect 14507 10965 14519 10999
rect 14461 10959 14519 10965
rect 14553 10999 14611 11005
rect 14553 10965 14565 10999
rect 14599 10996 14611 10999
rect 15010 10996 15016 11008
rect 14599 10968 15016 10996
rect 14599 10965 14611 10968
rect 14553 10959 14611 10965
rect 15010 10956 15016 10968
rect 15068 10956 15074 11008
rect 18230 10956 18236 11008
rect 18288 10996 18294 11008
rect 21634 10996 21640 11008
rect 18288 10968 21640 10996
rect 18288 10956 18294 10968
rect 21634 10956 21640 10968
rect 21692 10956 21698 11008
rect 25590 10956 25596 11008
rect 25648 10996 25654 11008
rect 26142 10996 26148 11008
rect 25648 10968 26148 10996
rect 25648 10956 25654 10968
rect 26142 10956 26148 10968
rect 26200 10996 26206 11008
rect 26528 10996 26556 11036
rect 26200 10968 26556 10996
rect 26200 10956 26206 10968
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 7558 10792 7564 10804
rect 7519 10764 7564 10792
rect 7558 10752 7564 10764
rect 7616 10752 7622 10804
rect 9677 10795 9735 10801
rect 9677 10761 9689 10795
rect 9723 10761 9735 10795
rect 9677 10755 9735 10761
rect 10413 10795 10471 10801
rect 10413 10761 10425 10795
rect 10459 10792 10471 10795
rect 11054 10792 11060 10804
rect 10459 10764 11060 10792
rect 10459 10761 10471 10764
rect 10413 10755 10471 10761
rect 8573 10727 8631 10733
rect 8573 10724 8585 10727
rect 7760 10696 8585 10724
rect 7760 10665 7788 10696
rect 8573 10693 8585 10696
rect 8619 10693 8631 10727
rect 8573 10687 8631 10693
rect 9217 10727 9275 10733
rect 9217 10693 9229 10727
rect 9263 10724 9275 10727
rect 9306 10724 9312 10736
rect 9263 10696 9312 10724
rect 9263 10693 9275 10696
rect 9217 10687 9275 10693
rect 9306 10684 9312 10696
rect 9364 10684 9370 10736
rect 9692 10724 9720 10755
rect 11054 10752 11060 10764
rect 11112 10752 11118 10804
rect 15378 10792 15384 10804
rect 12912 10764 15148 10792
rect 15339 10764 15384 10792
rect 12250 10724 12256 10736
rect 9692 10696 11928 10724
rect 7745 10659 7803 10665
rect 7745 10625 7757 10659
rect 7791 10625 7803 10659
rect 8202 10656 8208 10668
rect 8163 10628 8208 10656
rect 7745 10619 7803 10625
rect 8202 10616 8208 10628
rect 8260 10616 8266 10668
rect 8389 10659 8447 10665
rect 8389 10625 8401 10659
rect 8435 10625 8447 10659
rect 8389 10619 8447 10625
rect 8404 10452 8432 10619
rect 9122 10616 9128 10668
rect 9180 10656 9186 10668
rect 9493 10659 9551 10665
rect 9493 10656 9505 10659
rect 9180 10628 9505 10656
rect 9180 10616 9186 10628
rect 9493 10625 9505 10628
rect 9539 10625 9551 10659
rect 10778 10656 10784 10668
rect 10739 10628 10784 10656
rect 9493 10619 9551 10625
rect 10778 10616 10784 10628
rect 10836 10616 10842 10668
rect 11790 10656 11796 10668
rect 11751 10628 11796 10656
rect 11790 10616 11796 10628
rect 11848 10616 11854 10668
rect 11900 10665 11928 10696
rect 11992 10696 12256 10724
rect 11992 10665 12020 10696
rect 12250 10684 12256 10696
rect 12308 10684 12314 10736
rect 11885 10659 11943 10665
rect 11885 10625 11897 10659
rect 11931 10625 11943 10659
rect 11885 10619 11943 10625
rect 11977 10659 12035 10665
rect 11977 10625 11989 10659
rect 12023 10625 12035 10659
rect 11977 10619 12035 10625
rect 12158 10616 12164 10668
rect 12216 10656 12222 10668
rect 12912 10656 12940 10764
rect 14921 10727 14979 10733
rect 14921 10693 14933 10727
rect 14967 10724 14979 10727
rect 15010 10724 15016 10736
rect 14967 10696 15016 10724
rect 14967 10693 14979 10696
rect 14921 10687 14979 10693
rect 15010 10684 15016 10696
rect 15068 10684 15074 10736
rect 15120 10724 15148 10764
rect 15378 10752 15384 10764
rect 15436 10752 15442 10804
rect 15933 10795 15991 10801
rect 15933 10761 15945 10795
rect 15979 10792 15991 10795
rect 16114 10792 16120 10804
rect 15979 10764 16120 10792
rect 15979 10761 15991 10764
rect 15933 10755 15991 10761
rect 16114 10752 16120 10764
rect 16172 10752 16178 10804
rect 16850 10792 16856 10804
rect 16811 10764 16856 10792
rect 16850 10752 16856 10764
rect 16908 10752 16914 10804
rect 19797 10795 19855 10801
rect 19797 10792 19809 10795
rect 18064 10764 19809 10792
rect 17954 10724 17960 10736
rect 15120 10696 17960 10724
rect 17954 10684 17960 10696
rect 18012 10684 18018 10736
rect 18064 10733 18092 10764
rect 19797 10761 19809 10764
rect 19843 10761 19855 10795
rect 19797 10755 19855 10761
rect 19978 10752 19984 10804
rect 20036 10792 20042 10804
rect 20717 10795 20775 10801
rect 20717 10792 20729 10795
rect 20036 10764 20729 10792
rect 20036 10752 20042 10764
rect 20717 10761 20729 10764
rect 20763 10761 20775 10795
rect 20717 10755 20775 10761
rect 18049 10727 18107 10733
rect 18049 10693 18061 10727
rect 18095 10693 18107 10727
rect 18049 10687 18107 10693
rect 18141 10727 18199 10733
rect 18141 10693 18153 10727
rect 18187 10724 18199 10727
rect 18414 10724 18420 10736
rect 18187 10696 18420 10724
rect 18187 10693 18199 10696
rect 18141 10687 18199 10693
rect 18414 10684 18420 10696
rect 18472 10684 18478 10736
rect 19429 10727 19487 10733
rect 19429 10693 19441 10727
rect 19475 10693 19487 10727
rect 19429 10687 19487 10693
rect 19645 10727 19703 10733
rect 19645 10693 19657 10727
rect 19691 10724 19703 10727
rect 20257 10727 20315 10733
rect 20257 10724 20269 10727
rect 19691 10696 20269 10724
rect 19691 10693 19703 10696
rect 19645 10687 19703 10693
rect 20257 10693 20269 10696
rect 20303 10724 20315 10727
rect 20303 10696 22692 10724
rect 20303 10693 20315 10696
rect 20257 10687 20315 10693
rect 12216 10628 12940 10656
rect 13081 10659 13139 10665
rect 12216 10616 12222 10628
rect 13081 10625 13093 10659
rect 13127 10656 13139 10659
rect 13170 10656 13176 10668
rect 13127 10628 13176 10656
rect 13127 10625 13139 10628
rect 13081 10619 13139 10625
rect 13170 10616 13176 10628
rect 13228 10616 13234 10668
rect 13348 10659 13406 10665
rect 13348 10625 13360 10659
rect 13394 10656 13406 10659
rect 14826 10656 14832 10668
rect 13394 10628 14832 10656
rect 13394 10625 13406 10628
rect 13348 10619 13406 10625
rect 14826 10616 14832 10628
rect 14884 10616 14890 10668
rect 15197 10659 15255 10665
rect 15197 10625 15209 10659
rect 15243 10656 15255 10659
rect 15470 10656 15476 10668
rect 15243 10628 15476 10656
rect 15243 10625 15255 10628
rect 15197 10619 15255 10625
rect 15470 10616 15476 10628
rect 15528 10616 15534 10668
rect 15838 10656 15844 10668
rect 15799 10628 15844 10656
rect 15838 10616 15844 10628
rect 15896 10616 15902 10668
rect 17037 10659 17095 10665
rect 17037 10625 17049 10659
rect 17083 10656 17095 10659
rect 17773 10659 17831 10665
rect 17773 10656 17785 10659
rect 17083 10628 17785 10656
rect 17083 10625 17095 10628
rect 17037 10619 17095 10625
rect 17773 10625 17785 10628
rect 17819 10625 17831 10659
rect 17773 10619 17831 10625
rect 17974 10649 18032 10655
rect 17974 10615 17986 10649
rect 18020 10646 18032 10649
rect 18020 10618 18092 10646
rect 18020 10615 18032 10618
rect 17974 10609 18032 10615
rect 8478 10548 8484 10600
rect 8536 10588 8542 10600
rect 9309 10591 9367 10597
rect 9309 10588 9321 10591
rect 8536 10560 9321 10588
rect 8536 10548 8542 10560
rect 9309 10557 9321 10560
rect 9355 10557 9367 10591
rect 9309 10551 9367 10557
rect 10502 10548 10508 10600
rect 10560 10588 10566 10600
rect 10597 10591 10655 10597
rect 10597 10588 10609 10591
rect 10560 10560 10609 10588
rect 10560 10548 10566 10560
rect 10597 10557 10609 10560
rect 10643 10557 10655 10591
rect 10597 10551 10655 10557
rect 10686 10548 10692 10600
rect 10744 10588 10750 10600
rect 10873 10591 10931 10597
rect 10744 10560 10789 10588
rect 10744 10548 10750 10560
rect 10873 10557 10885 10591
rect 10919 10588 10931 10591
rect 11517 10591 11575 10597
rect 11517 10588 11529 10591
rect 10919 10560 11529 10588
rect 10919 10557 10931 10560
rect 10873 10551 10931 10557
rect 11517 10557 11529 10560
rect 11563 10557 11575 10591
rect 11517 10551 11575 10557
rect 14090 10548 14096 10600
rect 14148 10588 14154 10600
rect 14734 10588 14740 10600
rect 14148 10560 14740 10588
rect 14148 10548 14154 10560
rect 14734 10548 14740 10560
rect 14792 10588 14798 10600
rect 15013 10591 15071 10597
rect 15013 10588 15025 10591
rect 14792 10560 15025 10588
rect 14792 10548 14798 10560
rect 15013 10557 15025 10560
rect 15059 10557 15071 10591
rect 15013 10551 15071 10557
rect 17313 10591 17371 10597
rect 17313 10557 17325 10591
rect 17359 10557 17371 10591
rect 18064 10588 18092 10618
rect 18230 10616 18236 10668
rect 18288 10665 18294 10668
rect 18288 10659 18317 10665
rect 18305 10625 18317 10659
rect 19444 10656 19472 10687
rect 20162 10656 20168 10668
rect 19444 10628 20168 10656
rect 18288 10619 18317 10625
rect 18288 10616 18294 10619
rect 20162 10616 20168 10628
rect 20220 10616 20226 10668
rect 20533 10659 20591 10665
rect 20533 10625 20545 10659
rect 20579 10656 20591 10659
rect 21266 10656 21272 10668
rect 20579 10628 21272 10656
rect 20579 10625 20591 10628
rect 20533 10619 20591 10625
rect 21266 10616 21272 10628
rect 21324 10656 21330 10668
rect 21821 10659 21879 10665
rect 21821 10656 21833 10659
rect 21324 10628 21833 10656
rect 21324 10616 21330 10628
rect 21821 10625 21833 10628
rect 21867 10625 21879 10659
rect 21821 10619 21879 10625
rect 21910 10616 21916 10668
rect 21968 10656 21974 10668
rect 22005 10659 22063 10665
rect 22005 10656 22017 10659
rect 21968 10628 22017 10656
rect 21968 10616 21974 10628
rect 22005 10625 22017 10628
rect 22051 10625 22063 10659
rect 22005 10619 22063 10625
rect 18138 10588 18144 10600
rect 18064 10560 18144 10588
rect 17313 10551 17371 10557
rect 17328 10520 17356 10551
rect 18138 10548 18144 10560
rect 18196 10548 18202 10600
rect 18417 10591 18475 10597
rect 18417 10557 18429 10591
rect 18463 10588 18475 10591
rect 18506 10588 18512 10600
rect 18463 10560 18512 10588
rect 18463 10557 18475 10560
rect 18417 10551 18475 10557
rect 18506 10548 18512 10560
rect 18564 10548 18570 10600
rect 19886 10588 19892 10600
rect 18892 10560 19892 10588
rect 18892 10520 18920 10560
rect 19886 10548 19892 10560
rect 19944 10548 19950 10600
rect 20441 10591 20499 10597
rect 20441 10557 20453 10591
rect 20487 10588 20499 10591
rect 21358 10588 21364 10600
rect 20487 10560 21364 10588
rect 20487 10557 20499 10560
rect 20441 10551 20499 10557
rect 20456 10520 20484 10551
rect 21358 10548 21364 10560
rect 21416 10548 21422 10600
rect 17328 10492 18920 10520
rect 20088 10492 20484 10520
rect 22020 10520 22048 10619
rect 22664 10600 22692 10696
rect 23566 10684 23572 10736
rect 23624 10724 23630 10736
rect 24305 10727 24363 10733
rect 24305 10724 24317 10727
rect 23624 10696 24317 10724
rect 23624 10684 23630 10696
rect 24305 10693 24317 10696
rect 24351 10693 24363 10727
rect 24305 10687 24363 10693
rect 22833 10659 22891 10665
rect 22833 10625 22845 10659
rect 22879 10625 22891 10659
rect 22833 10619 22891 10625
rect 22646 10588 22652 10600
rect 22607 10560 22652 10588
rect 22646 10548 22652 10560
rect 22704 10548 22710 10600
rect 22848 10520 22876 10619
rect 25682 10616 25688 10668
rect 25740 10656 25746 10668
rect 26053 10659 26111 10665
rect 26053 10656 26065 10659
rect 25740 10628 26065 10656
rect 25740 10616 25746 10628
rect 26053 10625 26065 10628
rect 26099 10625 26111 10659
rect 26326 10656 26332 10668
rect 26287 10628 26332 10656
rect 26053 10619 26111 10625
rect 26326 10616 26332 10628
rect 26384 10616 26390 10668
rect 24765 10591 24823 10597
rect 24765 10557 24777 10591
rect 24811 10588 24823 10591
rect 26237 10591 26295 10597
rect 26237 10588 26249 10591
rect 24811 10560 26249 10588
rect 24811 10557 24823 10560
rect 24765 10551 24823 10557
rect 26237 10557 26249 10560
rect 26283 10588 26295 10591
rect 26510 10588 26516 10600
rect 26283 10560 26516 10588
rect 26283 10557 26295 10560
rect 26237 10551 26295 10557
rect 26510 10548 26516 10560
rect 26568 10548 26574 10600
rect 22020 10492 22876 10520
rect 9217 10455 9275 10461
rect 9217 10452 9229 10455
rect 8404 10424 9229 10452
rect 9217 10421 9229 10424
rect 9263 10452 9275 10455
rect 9306 10452 9312 10464
rect 9263 10424 9312 10452
rect 9263 10421 9275 10424
rect 9217 10415 9275 10421
rect 9306 10412 9312 10424
rect 9364 10412 9370 10464
rect 14182 10412 14188 10464
rect 14240 10452 14246 10464
rect 14366 10452 14372 10464
rect 14240 10424 14372 10452
rect 14240 10412 14246 10424
rect 14366 10412 14372 10424
rect 14424 10452 14430 10464
rect 14461 10455 14519 10461
rect 14461 10452 14473 10455
rect 14424 10424 14473 10452
rect 14424 10412 14430 10424
rect 14461 10421 14473 10424
rect 14507 10452 14519 10455
rect 14921 10455 14979 10461
rect 14921 10452 14933 10455
rect 14507 10424 14933 10452
rect 14507 10421 14519 10424
rect 14461 10415 14519 10421
rect 14921 10421 14933 10424
rect 14967 10421 14979 10455
rect 14921 10415 14979 10421
rect 17221 10455 17279 10461
rect 17221 10421 17233 10455
rect 17267 10452 17279 10455
rect 17954 10452 17960 10464
rect 17267 10424 17960 10452
rect 17267 10421 17279 10424
rect 17221 10415 17279 10421
rect 17954 10412 17960 10424
rect 18012 10412 18018 10464
rect 19613 10455 19671 10461
rect 19613 10421 19625 10455
rect 19659 10452 19671 10455
rect 20088 10452 20116 10492
rect 24210 10480 24216 10532
rect 24268 10520 24274 10532
rect 24581 10523 24639 10529
rect 24581 10520 24593 10523
rect 24268 10492 24593 10520
rect 24268 10480 24274 10492
rect 24581 10489 24593 10492
rect 24627 10489 24639 10523
rect 26142 10520 26148 10532
rect 26200 10529 26206 10532
rect 26107 10492 26148 10520
rect 24581 10483 24639 10489
rect 26142 10480 26148 10492
rect 26200 10483 26207 10529
rect 26200 10480 26206 10483
rect 19659 10424 20116 10452
rect 19659 10421 19671 10424
rect 19613 10415 19671 10421
rect 20162 10412 20168 10464
rect 20220 10452 20226 10464
rect 20257 10455 20315 10461
rect 20257 10452 20269 10455
rect 20220 10424 20269 10452
rect 20220 10412 20226 10424
rect 20257 10421 20269 10424
rect 20303 10421 20315 10455
rect 20257 10415 20315 10421
rect 22189 10455 22247 10461
rect 22189 10421 22201 10455
rect 22235 10452 22247 10455
rect 22278 10452 22284 10464
rect 22235 10424 22284 10452
rect 22235 10421 22247 10424
rect 22189 10415 22247 10421
rect 22278 10412 22284 10424
rect 22336 10412 22342 10464
rect 22922 10412 22928 10464
rect 22980 10452 22986 10464
rect 23017 10455 23075 10461
rect 23017 10452 23029 10455
rect 22980 10424 23029 10452
rect 22980 10412 22986 10424
rect 23017 10421 23029 10424
rect 23063 10421 23075 10455
rect 23017 10415 23075 10421
rect 25869 10455 25927 10461
rect 25869 10421 25881 10455
rect 25915 10452 25927 10455
rect 35802 10452 35808 10464
rect 25915 10424 35808 10452
rect 25915 10421 25927 10424
rect 25869 10415 25927 10421
rect 35802 10412 35808 10424
rect 35860 10412 35866 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 8389 10251 8447 10257
rect 8389 10217 8401 10251
rect 8435 10248 8447 10251
rect 8662 10248 8668 10260
rect 8435 10220 8668 10248
rect 8435 10217 8447 10220
rect 8389 10211 8447 10217
rect 8662 10208 8668 10220
rect 8720 10208 8726 10260
rect 10321 10251 10379 10257
rect 10321 10217 10333 10251
rect 10367 10217 10379 10251
rect 10502 10248 10508 10260
rect 10463 10220 10508 10248
rect 10321 10211 10379 10217
rect 8202 10140 8208 10192
rect 8260 10140 8266 10192
rect 8018 10112 8024 10124
rect 7931 10084 8024 10112
rect 8018 10072 8024 10084
rect 8076 10112 8082 10124
rect 8220 10112 8248 10140
rect 8076 10084 8248 10112
rect 10336 10112 10364 10211
rect 10502 10208 10508 10220
rect 10560 10208 10566 10260
rect 14826 10208 14832 10260
rect 14884 10248 14890 10260
rect 14921 10251 14979 10257
rect 14921 10248 14933 10251
rect 14884 10220 14933 10248
rect 14884 10208 14890 10220
rect 14921 10217 14933 10220
rect 14967 10217 14979 10251
rect 14921 10211 14979 10217
rect 16666 10208 16672 10260
rect 16724 10248 16730 10260
rect 17037 10251 17095 10257
rect 17037 10248 17049 10251
rect 16724 10220 17049 10248
rect 16724 10208 16730 10220
rect 17037 10217 17049 10220
rect 17083 10217 17095 10251
rect 17037 10211 17095 10217
rect 17773 10251 17831 10257
rect 17773 10217 17785 10251
rect 17819 10217 17831 10251
rect 17954 10248 17960 10260
rect 17915 10220 17960 10248
rect 17773 10211 17831 10217
rect 15102 10140 15108 10192
rect 15160 10180 15166 10192
rect 15160 10152 15700 10180
rect 15160 10140 15166 10152
rect 10336 10084 11100 10112
rect 8076 10072 8082 10084
rect 8205 10047 8263 10053
rect 8205 10013 8217 10047
rect 8251 10044 8263 10047
rect 8386 10044 8392 10056
rect 8251 10016 8392 10044
rect 8251 10013 8263 10016
rect 8205 10007 8263 10013
rect 8386 10004 8392 10016
rect 8444 10004 8450 10056
rect 9306 10044 9312 10056
rect 9267 10016 9312 10044
rect 9306 10004 9312 10016
rect 9364 10004 9370 10056
rect 9398 10004 9404 10056
rect 9456 10044 9462 10056
rect 9493 10047 9551 10053
rect 9493 10044 9505 10047
rect 9456 10016 9505 10044
rect 9456 10004 9462 10016
rect 9493 10013 9505 10016
rect 9539 10013 9551 10047
rect 9493 10007 9551 10013
rect 10318 10004 10324 10056
rect 10376 10044 10382 10056
rect 10870 10044 10876 10056
rect 10376 10016 10876 10044
rect 10376 10004 10382 10016
rect 10870 10004 10876 10016
rect 10928 10044 10934 10056
rect 10965 10047 11023 10053
rect 10965 10044 10977 10047
rect 10928 10016 10977 10044
rect 10928 10004 10934 10016
rect 10965 10013 10977 10016
rect 11011 10013 11023 10047
rect 11072 10044 11100 10084
rect 12250 10072 12256 10124
rect 12308 10112 12314 10124
rect 15194 10112 15200 10124
rect 12308 10084 13032 10112
rect 12308 10072 12314 10084
rect 11606 10044 11612 10056
rect 11072 10016 11612 10044
rect 10965 10007 11023 10013
rect 11606 10004 11612 10016
rect 11664 10004 11670 10056
rect 12894 10044 12900 10056
rect 12855 10016 12900 10044
rect 12894 10004 12900 10016
rect 12952 10004 12958 10056
rect 13004 10053 13032 10084
rect 14292 10084 15200 10112
rect 12989 10047 13047 10053
rect 12989 10013 13001 10047
rect 13035 10013 13047 10047
rect 14182 10044 14188 10056
rect 14143 10016 14188 10044
rect 12989 10007 13047 10013
rect 14182 10004 14188 10016
rect 14240 10004 14246 10056
rect 14292 10053 14320 10084
rect 15194 10072 15200 10084
rect 15252 10072 15258 10124
rect 15672 10121 15700 10152
rect 15657 10115 15715 10121
rect 15657 10081 15669 10115
rect 15703 10081 15715 10115
rect 15657 10075 15715 10081
rect 14277 10047 14335 10053
rect 14277 10013 14289 10047
rect 14323 10013 14335 10047
rect 14277 10007 14335 10013
rect 14366 10004 14372 10056
rect 14424 10044 14430 10056
rect 15105 10047 15163 10053
rect 15105 10044 15117 10047
rect 14424 10016 15117 10044
rect 14424 10004 14430 10016
rect 15105 10013 15117 10016
rect 15151 10013 15163 10047
rect 15672 10044 15700 10075
rect 17052 10044 17080 10211
rect 17788 10180 17816 10211
rect 17954 10208 17960 10220
rect 18012 10208 18018 10260
rect 20162 10208 20168 10260
rect 20220 10248 20226 10260
rect 20625 10251 20683 10257
rect 20625 10248 20637 10251
rect 20220 10220 20637 10248
rect 20220 10208 20226 10220
rect 20625 10217 20637 10220
rect 20671 10217 20683 10251
rect 20625 10211 20683 10217
rect 22646 10208 22652 10260
rect 22704 10248 22710 10260
rect 23017 10251 23075 10257
rect 23017 10248 23029 10251
rect 22704 10220 23029 10248
rect 22704 10208 22710 10220
rect 23017 10217 23029 10220
rect 23063 10217 23075 10251
rect 24578 10248 24584 10260
rect 24539 10220 24584 10248
rect 23017 10211 23075 10217
rect 24578 10208 24584 10220
rect 24636 10208 24642 10260
rect 25406 10248 25412 10260
rect 25367 10220 25412 10248
rect 25406 10208 25412 10220
rect 25464 10208 25470 10260
rect 18046 10180 18052 10192
rect 17788 10152 18052 10180
rect 18046 10140 18052 10152
rect 18104 10140 18110 10192
rect 24118 10140 24124 10192
rect 24176 10180 24182 10192
rect 24489 10183 24547 10189
rect 24489 10180 24501 10183
rect 24176 10152 24501 10180
rect 24176 10140 24182 10152
rect 24489 10149 24501 10152
rect 24535 10149 24547 10183
rect 24489 10143 24547 10149
rect 17681 10115 17739 10121
rect 17681 10081 17693 10115
rect 17727 10112 17739 10115
rect 19058 10112 19064 10124
rect 17727 10084 19064 10112
rect 17727 10081 17739 10084
rect 17681 10075 17739 10081
rect 19058 10072 19064 10084
rect 19116 10072 19122 10124
rect 20714 10072 20720 10124
rect 20772 10112 20778 10124
rect 21637 10115 21695 10121
rect 21637 10112 21649 10115
rect 20772 10084 21649 10112
rect 20772 10072 20778 10084
rect 21637 10081 21649 10084
rect 21683 10081 21695 10115
rect 24670 10112 24676 10124
rect 24631 10084 24676 10112
rect 21637 10075 21695 10081
rect 24670 10072 24676 10084
rect 24728 10072 24734 10124
rect 25590 10112 25596 10124
rect 25148 10084 25596 10112
rect 17497 10047 17555 10053
rect 17497 10044 17509 10047
rect 15672 10016 16620 10044
rect 17052 10016 17509 10044
rect 15105 10007 15163 10013
rect 8404 9908 8432 10004
rect 16592 9988 16620 10016
rect 17497 10013 17509 10016
rect 17543 10013 17555 10047
rect 17770 10044 17776 10056
rect 17731 10016 17776 10044
rect 17497 10007 17555 10013
rect 17770 10004 17776 10016
rect 17828 10004 17834 10056
rect 18598 10044 18604 10056
rect 18559 10016 18604 10044
rect 18598 10004 18604 10016
rect 18656 10004 18662 10056
rect 19242 10044 19248 10056
rect 19203 10016 19248 10044
rect 19242 10004 19248 10016
rect 19300 10004 19306 10056
rect 19334 10004 19340 10056
rect 19392 10044 19398 10056
rect 19501 10047 19559 10053
rect 19501 10044 19513 10047
rect 19392 10016 19513 10044
rect 19392 10004 19398 10016
rect 19501 10013 19513 10016
rect 19547 10013 19559 10047
rect 19501 10007 19559 10013
rect 24397 10047 24455 10053
rect 24397 10013 24409 10047
rect 24443 10044 24455 10047
rect 25148 10044 25176 10084
rect 25590 10072 25596 10084
rect 25648 10072 25654 10124
rect 25314 10044 25320 10056
rect 24443 10016 25176 10044
rect 25275 10016 25320 10044
rect 24443 10013 24455 10016
rect 24397 10007 24455 10013
rect 25314 10004 25320 10016
rect 25372 10004 25378 10056
rect 25501 10047 25559 10053
rect 25501 10013 25513 10047
rect 25547 10044 25559 10047
rect 25682 10044 25688 10056
rect 25547 10016 25688 10044
rect 25547 10013 25559 10016
rect 25501 10007 25559 10013
rect 25682 10004 25688 10016
rect 25740 10004 25746 10056
rect 9122 9976 9128 9988
rect 9083 9948 9128 9976
rect 9122 9936 9128 9948
rect 9180 9936 9186 9988
rect 10137 9979 10195 9985
rect 10137 9945 10149 9979
rect 10183 9976 10195 9979
rect 10183 9948 10640 9976
rect 10183 9945 10195 9948
rect 10137 9939 10195 9945
rect 9401 9911 9459 9917
rect 9401 9908 9413 9911
rect 8404 9880 9413 9908
rect 9401 9877 9413 9880
rect 9447 9877 9459 9911
rect 9401 9871 9459 9877
rect 9677 9911 9735 9917
rect 9677 9877 9689 9911
rect 9723 9908 9735 9911
rect 10337 9911 10395 9917
rect 10337 9908 10349 9911
rect 9723 9880 10349 9908
rect 9723 9877 9735 9880
rect 9677 9871 9735 9877
rect 10337 9877 10349 9880
rect 10383 9877 10395 9911
rect 10612 9908 10640 9948
rect 10686 9936 10692 9988
rect 10744 9976 10750 9988
rect 11210 9979 11268 9985
rect 11210 9976 11222 9979
rect 10744 9948 11222 9976
rect 10744 9936 10750 9948
rect 11210 9945 11222 9948
rect 11256 9945 11268 9979
rect 11210 9939 11268 9945
rect 11330 9936 11336 9988
rect 11388 9976 11394 9988
rect 13173 9979 13231 9985
rect 13173 9976 13185 9979
rect 11388 9948 13185 9976
rect 11388 9936 11394 9948
rect 13173 9945 13185 9948
rect 13219 9945 13231 9979
rect 13173 9939 13231 9945
rect 14461 9979 14519 9985
rect 14461 9945 14473 9979
rect 14507 9976 14519 9979
rect 15378 9976 15384 9988
rect 14507 9948 15384 9976
rect 14507 9945 14519 9948
rect 14461 9939 14519 9945
rect 15378 9936 15384 9948
rect 15436 9936 15442 9988
rect 15930 9985 15936 9988
rect 15924 9939 15936 9985
rect 15988 9976 15994 9988
rect 15988 9948 16024 9976
rect 15930 9936 15936 9939
rect 15988 9936 15994 9948
rect 16574 9936 16580 9988
rect 16632 9936 16638 9988
rect 21904 9979 21962 9985
rect 21904 9945 21916 9979
rect 21950 9976 21962 9979
rect 22094 9976 22100 9988
rect 21950 9948 22100 9976
rect 21950 9945 21962 9948
rect 21904 9939 21962 9945
rect 22094 9936 22100 9948
rect 22152 9936 22158 9988
rect 11514 9908 11520 9920
rect 10612 9880 11520 9908
rect 10337 9871 10395 9877
rect 11514 9868 11520 9880
rect 11572 9908 11578 9920
rect 12342 9908 12348 9920
rect 11572 9880 12348 9908
rect 11572 9868 11578 9880
rect 12342 9868 12348 9880
rect 12400 9868 12406 9920
rect 18414 9908 18420 9920
rect 18375 9880 18420 9908
rect 18414 9868 18420 9880
rect 18472 9868 18478 9920
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 8573 9707 8631 9713
rect 8573 9673 8585 9707
rect 8619 9704 8631 9707
rect 9306 9704 9312 9716
rect 8619 9676 9312 9704
rect 8619 9673 8631 9676
rect 8573 9667 8631 9673
rect 9306 9664 9312 9676
rect 9364 9664 9370 9716
rect 10686 9664 10692 9716
rect 10744 9704 10750 9716
rect 10781 9707 10839 9713
rect 10781 9704 10793 9707
rect 10744 9676 10793 9704
rect 10744 9664 10750 9676
rect 10781 9673 10793 9676
rect 10827 9673 10839 9707
rect 10781 9667 10839 9673
rect 11790 9664 11796 9716
rect 11848 9704 11854 9716
rect 11977 9707 12035 9713
rect 11977 9704 11989 9707
rect 11848 9676 11989 9704
rect 11848 9664 11854 9676
rect 11977 9673 11989 9676
rect 12023 9673 12035 9707
rect 15930 9704 15936 9716
rect 15891 9676 15936 9704
rect 11977 9667 12035 9673
rect 15930 9664 15936 9676
rect 15988 9664 15994 9716
rect 17696 9676 19288 9704
rect 10318 9636 10324 9648
rect 7208 9608 10324 9636
rect 7208 9577 7236 9608
rect 10318 9596 10324 9608
rect 10376 9596 10382 9648
rect 10870 9596 10876 9648
rect 10928 9636 10934 9648
rect 11517 9639 11575 9645
rect 11517 9636 11529 9639
rect 10928 9608 11529 9636
rect 10928 9596 10934 9608
rect 11517 9605 11529 9608
rect 11563 9605 11575 9639
rect 17037 9639 17095 9645
rect 17037 9636 17049 9639
rect 11517 9599 11575 9605
rect 16132 9608 17049 9636
rect 7193 9571 7251 9577
rect 7193 9537 7205 9571
rect 7239 9537 7251 9571
rect 7193 9531 7251 9537
rect 7460 9571 7518 9577
rect 7460 9537 7472 9571
rect 7506 9568 7518 9571
rect 9214 9568 9220 9580
rect 7506 9540 9076 9568
rect 9175 9540 9220 9568
rect 7506 9537 7518 9540
rect 7460 9531 7518 9537
rect 9048 9441 9076 9540
rect 9214 9528 9220 9540
rect 9272 9528 9278 9580
rect 10965 9571 11023 9577
rect 10965 9537 10977 9571
rect 11011 9568 11023 9571
rect 11330 9568 11336 9580
rect 11011 9540 11336 9568
rect 11011 9537 11023 9540
rect 10965 9531 11023 9537
rect 11330 9528 11336 9540
rect 11388 9528 11394 9580
rect 11422 9528 11428 9580
rect 11480 9568 11486 9580
rect 11793 9571 11851 9577
rect 11793 9568 11805 9571
rect 11480 9540 11805 9568
rect 11480 9528 11486 9540
rect 11793 9537 11805 9540
rect 11839 9568 11851 9571
rect 12250 9568 12256 9580
rect 11839 9540 12256 9568
rect 11839 9537 11851 9540
rect 11793 9531 11851 9537
rect 12250 9528 12256 9540
rect 12308 9528 12314 9580
rect 13078 9528 13084 9580
rect 13136 9568 13142 9580
rect 13357 9571 13415 9577
rect 13357 9568 13369 9571
rect 13136 9540 13369 9568
rect 13136 9528 13142 9540
rect 13357 9537 13369 9540
rect 13403 9537 13415 9571
rect 13357 9531 13415 9537
rect 13624 9571 13682 9577
rect 13624 9537 13636 9571
rect 13670 9568 13682 9571
rect 15378 9568 15384 9580
rect 13670 9540 15240 9568
rect 15339 9540 15384 9568
rect 13670 9537 13682 9540
rect 13624 9531 13682 9537
rect 11606 9500 11612 9512
rect 11567 9472 11612 9500
rect 11606 9460 11612 9472
rect 11664 9460 11670 9512
rect 15212 9441 15240 9540
rect 15378 9528 15384 9540
rect 15436 9528 15442 9580
rect 16132 9577 16160 9608
rect 17037 9605 17049 9608
rect 17083 9605 17095 9639
rect 17037 9599 17095 9605
rect 17696 9577 17724 9676
rect 19260 9648 19288 9676
rect 17948 9639 18006 9645
rect 17948 9605 17960 9639
rect 17994 9636 18006 9639
rect 18414 9636 18420 9648
rect 17994 9608 18420 9636
rect 17994 9605 18006 9608
rect 17948 9599 18006 9605
rect 18414 9596 18420 9608
rect 18472 9596 18478 9648
rect 19242 9596 19248 9648
rect 19300 9636 19306 9648
rect 20714 9636 20720 9648
rect 19300 9608 20720 9636
rect 19300 9596 19306 9608
rect 19904 9577 19932 9608
rect 20714 9596 20720 9608
rect 20772 9636 20778 9648
rect 20772 9608 22232 9636
rect 20772 9596 20778 9608
rect 16117 9571 16175 9577
rect 16117 9537 16129 9571
rect 16163 9537 16175 9571
rect 16853 9571 16911 9577
rect 16853 9568 16865 9571
rect 16117 9531 16175 9537
rect 16546 9540 16865 9568
rect 15286 9460 15292 9512
rect 15344 9500 15350 9512
rect 16206 9500 16212 9512
rect 15344 9472 16212 9500
rect 15344 9460 15350 9472
rect 16206 9460 16212 9472
rect 16264 9500 16270 9512
rect 16546 9500 16574 9540
rect 16853 9537 16865 9540
rect 16899 9537 16911 9571
rect 16853 9531 16911 9537
rect 17681 9571 17739 9577
rect 17681 9537 17693 9571
rect 17727 9537 17739 9571
rect 17681 9531 17739 9537
rect 19889 9571 19947 9577
rect 19889 9537 19901 9571
rect 19935 9537 19947 9571
rect 19889 9531 19947 9537
rect 20156 9571 20214 9577
rect 20156 9537 20168 9571
rect 20202 9568 20214 9571
rect 20990 9568 20996 9580
rect 20202 9540 20996 9568
rect 20202 9537 20214 9540
rect 20156 9531 20214 9537
rect 20990 9528 20996 9540
rect 21048 9528 21054 9580
rect 22204 9577 22232 9608
rect 22189 9571 22247 9577
rect 22189 9537 22201 9571
rect 22235 9537 22247 9571
rect 22189 9531 22247 9537
rect 22456 9571 22514 9577
rect 22456 9537 22468 9571
rect 22502 9568 22514 9571
rect 22738 9568 22744 9580
rect 22502 9540 22744 9568
rect 22502 9537 22514 9540
rect 22456 9531 22514 9537
rect 22738 9528 22744 9540
rect 22796 9528 22802 9580
rect 16666 9500 16672 9512
rect 16264 9472 16574 9500
rect 16627 9472 16672 9500
rect 16264 9460 16270 9472
rect 16666 9460 16672 9472
rect 16724 9460 16730 9512
rect 9033 9435 9091 9441
rect 9033 9401 9045 9435
rect 9079 9401 9091 9435
rect 9033 9395 9091 9401
rect 15197 9435 15255 9441
rect 15197 9401 15209 9435
rect 15243 9401 15255 9435
rect 19058 9432 19064 9444
rect 19019 9404 19064 9432
rect 15197 9395 15255 9401
rect 19058 9392 19064 9404
rect 19116 9392 19122 9444
rect 11514 9364 11520 9376
rect 11475 9336 11520 9364
rect 11514 9324 11520 9336
rect 11572 9324 11578 9376
rect 14734 9364 14740 9376
rect 14695 9336 14740 9364
rect 14734 9324 14740 9336
rect 14792 9324 14798 9376
rect 21266 9364 21272 9376
rect 21227 9336 21272 9364
rect 21266 9324 21272 9336
rect 21324 9324 21330 9376
rect 21358 9324 21364 9376
rect 21416 9364 21422 9376
rect 23569 9367 23627 9373
rect 23569 9364 23581 9367
rect 21416 9336 23581 9364
rect 21416 9324 21422 9336
rect 23569 9333 23581 9336
rect 23615 9333 23627 9367
rect 23569 9327 23627 9333
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 8389 9163 8447 9169
rect 8389 9129 8401 9163
rect 8435 9160 8447 9163
rect 9214 9160 9220 9172
rect 8435 9132 9220 9160
rect 8435 9129 8447 9132
rect 8389 9123 8447 9129
rect 9214 9120 9220 9132
rect 9272 9120 9278 9172
rect 15010 9120 15016 9172
rect 15068 9160 15074 9172
rect 15473 9163 15531 9169
rect 15473 9160 15485 9163
rect 15068 9132 15485 9160
rect 15068 9120 15074 9132
rect 15473 9129 15485 9132
rect 15519 9129 15531 9163
rect 15473 9123 15531 9129
rect 18138 9120 18144 9172
rect 18196 9160 18202 9172
rect 18601 9163 18659 9169
rect 18601 9160 18613 9163
rect 18196 9132 18613 9160
rect 18196 9120 18202 9132
rect 18601 9129 18613 9132
rect 18647 9129 18659 9163
rect 18601 9123 18659 9129
rect 19426 9120 19432 9172
rect 19484 9160 19490 9172
rect 19613 9163 19671 9169
rect 19613 9160 19625 9163
rect 19484 9132 19625 9160
rect 19484 9120 19490 9132
rect 19613 9129 19625 9132
rect 19659 9129 19671 9163
rect 20990 9160 20996 9172
rect 20951 9132 20996 9160
rect 19613 9123 19671 9129
rect 20990 9120 20996 9132
rect 21048 9120 21054 9172
rect 22094 9160 22100 9172
rect 22055 9132 22100 9160
rect 22094 9120 22100 9132
rect 22152 9120 22158 9172
rect 22738 9160 22744 9172
rect 22699 9132 22744 9160
rect 22738 9120 22744 9132
rect 22796 9120 22802 9172
rect 16666 9052 16672 9104
rect 16724 9092 16730 9104
rect 17770 9092 17776 9104
rect 16724 9064 17776 9092
rect 16724 9052 16730 9064
rect 17770 9052 17776 9064
rect 17828 9092 17834 9104
rect 18049 9095 18107 9101
rect 18049 9092 18061 9095
rect 17828 9064 18061 9092
rect 17828 9052 17834 9064
rect 18049 9061 18061 9064
rect 18095 9061 18107 9095
rect 18049 9055 18107 9061
rect 8018 9024 8024 9036
rect 7979 8996 8024 9024
rect 8018 8984 8024 8996
rect 8076 9024 8082 9036
rect 9493 9027 9551 9033
rect 9493 9024 9505 9027
rect 8076 8996 9505 9024
rect 8076 8984 8082 8996
rect 9493 8993 9505 8996
rect 9539 8993 9551 9027
rect 9493 8987 9551 8993
rect 12161 9027 12219 9033
rect 12161 8993 12173 9027
rect 12207 9024 12219 9027
rect 12250 9024 12256 9036
rect 12207 8996 12256 9024
rect 12207 8993 12219 8996
rect 12161 8987 12219 8993
rect 12250 8984 12256 8996
rect 12308 8984 12314 9036
rect 20162 9024 20168 9036
rect 20123 8996 20168 9024
rect 20162 8984 20168 8996
rect 20220 8984 20226 9036
rect 21910 9024 21916 9036
rect 20364 8996 21916 9024
rect 8205 8959 8263 8965
rect 8205 8925 8217 8959
rect 8251 8956 8263 8959
rect 8294 8956 8300 8968
rect 8251 8928 8300 8956
rect 8251 8925 8263 8928
rect 8205 8919 8263 8925
rect 8294 8916 8300 8928
rect 8352 8916 8358 8968
rect 9677 8959 9735 8965
rect 9677 8925 9689 8959
rect 9723 8925 9735 8959
rect 10318 8956 10324 8968
rect 10279 8928 10324 8956
rect 9677 8919 9735 8925
rect 9692 8888 9720 8919
rect 10318 8916 10324 8928
rect 10376 8916 10382 8968
rect 12342 8956 12348 8968
rect 12303 8928 12348 8956
rect 12342 8916 12348 8928
rect 12400 8916 12406 8968
rect 13538 8956 13544 8968
rect 13499 8928 13544 8956
rect 13538 8916 13544 8928
rect 13596 8916 13602 8968
rect 13722 8916 13728 8968
rect 13780 8956 13786 8968
rect 14093 8959 14151 8965
rect 14093 8956 14105 8959
rect 13780 8928 14105 8956
rect 13780 8916 13786 8928
rect 14093 8925 14105 8928
rect 14139 8925 14151 8959
rect 14093 8919 14151 8925
rect 16025 8959 16083 8965
rect 16025 8925 16037 8959
rect 16071 8925 16083 8959
rect 16025 8919 16083 8925
rect 16117 8959 16175 8965
rect 16117 8925 16129 8959
rect 16163 8956 16175 8959
rect 16206 8956 16212 8968
rect 16163 8928 16212 8956
rect 16163 8925 16175 8928
rect 16117 8919 16175 8925
rect 10588 8891 10646 8897
rect 9692 8860 10548 8888
rect 9861 8823 9919 8829
rect 9861 8789 9873 8823
rect 9907 8820 9919 8823
rect 10226 8820 10232 8832
rect 9907 8792 10232 8820
rect 9907 8789 9919 8792
rect 9861 8783 9919 8789
rect 10226 8780 10232 8792
rect 10284 8780 10290 8832
rect 10520 8820 10548 8860
rect 10588 8857 10600 8891
rect 10634 8888 10646 8891
rect 10686 8888 10692 8900
rect 10634 8860 10692 8888
rect 10634 8857 10646 8860
rect 10588 8851 10646 8857
rect 10686 8848 10692 8860
rect 10744 8848 10750 8900
rect 14338 8891 14396 8897
rect 14338 8888 14350 8891
rect 13372 8860 14350 8888
rect 10870 8820 10876 8832
rect 10520 8792 10876 8820
rect 10870 8780 10876 8792
rect 10928 8820 10934 8832
rect 11701 8823 11759 8829
rect 11701 8820 11713 8823
rect 10928 8792 11713 8820
rect 10928 8780 10934 8792
rect 11701 8789 11713 8792
rect 11747 8789 11759 8823
rect 12526 8820 12532 8832
rect 12487 8792 12532 8820
rect 11701 8783 11759 8789
rect 12526 8780 12532 8792
rect 12584 8780 12590 8832
rect 13372 8829 13400 8860
rect 14338 8857 14350 8860
rect 14384 8857 14396 8891
rect 16040 8888 16068 8919
rect 16206 8916 16212 8928
rect 16264 8916 16270 8968
rect 16301 8959 16359 8965
rect 16301 8925 16313 8959
rect 16347 8956 16359 8959
rect 16945 8959 17003 8965
rect 16945 8956 16957 8959
rect 16347 8928 16957 8956
rect 16347 8925 16359 8928
rect 16301 8919 16359 8925
rect 16945 8925 16957 8928
rect 16991 8925 17003 8959
rect 16945 8919 17003 8925
rect 18325 8959 18383 8965
rect 18325 8925 18337 8959
rect 18371 8956 18383 8959
rect 19058 8956 19064 8968
rect 18371 8928 19064 8956
rect 18371 8925 18383 8928
rect 18325 8919 18383 8925
rect 19058 8916 19064 8928
rect 19116 8956 19122 8968
rect 20364 8965 20392 8996
rect 21910 8984 21916 8996
rect 21968 8984 21974 9036
rect 19245 8959 19303 8965
rect 19245 8956 19257 8959
rect 19116 8928 19257 8956
rect 19116 8916 19122 8928
rect 19245 8925 19257 8928
rect 19291 8925 19303 8959
rect 19245 8919 19303 8925
rect 19429 8959 19487 8965
rect 19429 8925 19441 8959
rect 19475 8956 19487 8959
rect 20349 8959 20407 8965
rect 20349 8956 20361 8959
rect 19475 8928 20361 8956
rect 19475 8925 19487 8928
rect 19429 8919 19487 8925
rect 20349 8925 20361 8928
rect 20395 8925 20407 8959
rect 20349 8919 20407 8925
rect 20533 8959 20591 8965
rect 20533 8925 20545 8959
rect 20579 8956 20591 8959
rect 21177 8959 21235 8965
rect 21177 8956 21189 8959
rect 20579 8928 21189 8956
rect 20579 8925 20591 8928
rect 20533 8919 20591 8925
rect 21177 8925 21189 8928
rect 21223 8925 21235 8959
rect 22278 8956 22284 8968
rect 22239 8928 22284 8956
rect 21177 8919 21235 8925
rect 22278 8916 22284 8928
rect 22336 8916 22342 8968
rect 22922 8956 22928 8968
rect 22883 8928 22928 8956
rect 22922 8916 22928 8928
rect 22980 8916 22986 8968
rect 18046 8888 18052 8900
rect 16040 8860 18052 8888
rect 14338 8851 14396 8857
rect 18046 8848 18052 8860
rect 18104 8888 18110 8900
rect 18417 8891 18475 8897
rect 18104 8860 18276 8888
rect 18104 8848 18110 8860
rect 13357 8823 13415 8829
rect 13357 8789 13369 8823
rect 13403 8789 13415 8823
rect 16758 8820 16764 8832
rect 16719 8792 16764 8820
rect 13357 8783 13415 8789
rect 16758 8780 16764 8792
rect 16816 8780 16822 8832
rect 18248 8829 18276 8860
rect 18417 8857 18429 8891
rect 18463 8888 18475 8891
rect 21266 8888 21272 8900
rect 18463 8860 21272 8888
rect 18463 8857 18475 8860
rect 18417 8851 18475 8857
rect 21266 8848 21272 8860
rect 21324 8848 21330 8900
rect 18233 8823 18291 8829
rect 18233 8789 18245 8823
rect 18279 8820 18291 8823
rect 18598 8820 18604 8832
rect 18279 8792 18604 8820
rect 18279 8789 18291 8792
rect 18233 8783 18291 8789
rect 18598 8780 18604 8792
rect 18656 8780 18662 8832
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 8294 8576 8300 8628
rect 8352 8616 8358 8628
rect 9122 8616 9128 8628
rect 8352 8588 9128 8616
rect 8352 8576 8358 8588
rect 9122 8576 9128 8588
rect 9180 8616 9186 8628
rect 9585 8619 9643 8625
rect 9585 8616 9597 8619
rect 9180 8588 9597 8616
rect 9180 8576 9186 8588
rect 9585 8585 9597 8588
rect 9631 8585 9643 8619
rect 9585 8579 9643 8585
rect 10045 8619 10103 8625
rect 10045 8585 10057 8619
rect 10091 8585 10103 8619
rect 10686 8616 10692 8628
rect 10647 8588 10692 8616
rect 10045 8579 10103 8585
rect 8472 8551 8530 8557
rect 8472 8517 8484 8551
rect 8518 8548 8530 8551
rect 10060 8548 10088 8579
rect 10686 8576 10692 8588
rect 10744 8576 10750 8628
rect 11514 8576 11520 8628
rect 11572 8616 11578 8628
rect 13081 8619 13139 8625
rect 13081 8616 13093 8619
rect 11572 8588 13093 8616
rect 11572 8576 11578 8588
rect 13081 8585 13093 8588
rect 13127 8585 13139 8619
rect 13081 8579 13139 8585
rect 13538 8576 13544 8628
rect 13596 8616 13602 8628
rect 14185 8619 14243 8625
rect 14185 8616 14197 8619
rect 13596 8588 14197 8616
rect 13596 8576 13602 8588
rect 14185 8585 14197 8588
rect 14231 8585 14243 8619
rect 14185 8579 14243 8585
rect 16117 8619 16175 8625
rect 16117 8585 16129 8619
rect 16163 8616 16175 8619
rect 16666 8616 16672 8628
rect 16163 8588 16672 8616
rect 16163 8585 16175 8588
rect 16117 8579 16175 8585
rect 16666 8576 16672 8588
rect 16724 8576 16730 8628
rect 8518 8520 10088 8548
rect 8518 8517 8530 8520
rect 8472 8511 8530 8517
rect 10318 8508 10324 8560
rect 10376 8548 10382 8560
rect 13722 8548 13728 8560
rect 10376 8520 13728 8548
rect 10376 8508 10382 8520
rect 8205 8483 8263 8489
rect 8205 8449 8217 8483
rect 8251 8480 8263 8483
rect 10226 8480 10232 8492
rect 8251 8452 9812 8480
rect 10187 8452 10232 8480
rect 8251 8449 8263 8452
rect 8205 8443 8263 8449
rect 9784 8412 9812 8452
rect 10226 8440 10232 8452
rect 10284 8440 10290 8492
rect 10873 8483 10931 8489
rect 10873 8449 10885 8483
rect 10919 8480 10931 8483
rect 11606 8480 11612 8492
rect 10919 8452 11612 8480
rect 10919 8449 10931 8452
rect 10873 8443 10931 8449
rect 11606 8440 11612 8452
rect 11664 8440 11670 8492
rect 11716 8489 11744 8520
rect 13722 8508 13728 8520
rect 13780 8508 13786 8560
rect 14734 8548 14740 8560
rect 13924 8520 14740 8548
rect 11974 8489 11980 8492
rect 11701 8483 11759 8489
rect 11701 8449 11713 8483
rect 11747 8449 11759 8483
rect 11701 8443 11759 8449
rect 11968 8443 11980 8489
rect 12032 8480 12038 8492
rect 13924 8489 13952 8520
rect 14734 8508 14740 8520
rect 14792 8508 14798 8560
rect 15004 8551 15062 8557
rect 15004 8517 15016 8551
rect 15050 8548 15062 8551
rect 16758 8548 16764 8560
rect 15050 8520 16764 8548
rect 15050 8517 15062 8520
rect 15004 8511 15062 8517
rect 16758 8508 16764 8520
rect 16816 8508 16822 8560
rect 13909 8483 13967 8489
rect 12032 8452 12068 8480
rect 11974 8440 11980 8443
rect 12032 8440 12038 8452
rect 13909 8449 13921 8483
rect 13955 8449 13967 8483
rect 13909 8443 13967 8449
rect 14001 8483 14059 8489
rect 14001 8449 14013 8483
rect 14047 8480 14059 8483
rect 15286 8480 15292 8492
rect 14047 8452 15292 8480
rect 14047 8449 14059 8452
rect 14001 8443 14059 8449
rect 15286 8440 15292 8452
rect 15344 8440 15350 8492
rect 17313 8483 17371 8489
rect 17313 8449 17325 8483
rect 17359 8480 17371 8483
rect 17586 8480 17592 8492
rect 17359 8452 17592 8480
rect 17359 8449 17371 8452
rect 17313 8443 17371 8449
rect 17586 8440 17592 8452
rect 17644 8440 17650 8492
rect 10318 8412 10324 8424
rect 9784 8384 10324 8412
rect 10318 8372 10324 8384
rect 10376 8372 10382 8424
rect 13722 8372 13728 8424
rect 13780 8412 13786 8424
rect 14737 8415 14795 8421
rect 14737 8412 14749 8415
rect 13780 8384 14749 8412
rect 13780 8372 13786 8384
rect 14737 8381 14749 8384
rect 14783 8381 14795 8415
rect 14737 8375 14795 8381
rect 14752 8276 14780 8375
rect 16574 8344 16580 8356
rect 15672 8316 16580 8344
rect 15672 8276 15700 8316
rect 16574 8304 16580 8316
rect 16632 8304 16638 8356
rect 14752 8248 15700 8276
rect 17129 8279 17187 8285
rect 17129 8245 17141 8279
rect 17175 8276 17187 8279
rect 17310 8276 17316 8288
rect 17175 8248 17316 8276
rect 17175 8245 17187 8248
rect 17129 8239 17187 8245
rect 17310 8236 17316 8248
rect 17368 8236 17374 8288
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 10873 8075 10931 8081
rect 10873 8041 10885 8075
rect 10919 8072 10931 8075
rect 11422 8072 11428 8084
rect 10919 8044 11428 8072
rect 10919 8041 10931 8044
rect 10873 8035 10931 8041
rect 11422 8032 11428 8044
rect 11480 8032 11486 8084
rect 11606 8032 11612 8084
rect 11664 8072 11670 8084
rect 11701 8075 11759 8081
rect 11701 8072 11713 8075
rect 11664 8044 11713 8072
rect 11664 8032 11670 8044
rect 11701 8041 11713 8044
rect 11747 8041 11759 8075
rect 11701 8035 11759 8041
rect 11974 8032 11980 8084
rect 12032 8072 12038 8084
rect 12161 8075 12219 8081
rect 12161 8072 12173 8075
rect 12032 8044 12173 8072
rect 12032 8032 12038 8044
rect 12161 8041 12173 8044
rect 12207 8041 12219 8075
rect 12161 8035 12219 8041
rect 12250 8032 12256 8084
rect 12308 8072 12314 8084
rect 17218 8072 17224 8084
rect 12308 8044 17224 8072
rect 12308 8032 12314 8044
rect 17218 8032 17224 8044
rect 17276 8032 17282 8084
rect 18598 8072 18604 8084
rect 18559 8044 18604 8072
rect 18598 8032 18604 8044
rect 18656 8032 18662 8084
rect 11330 7936 11336 7948
rect 11243 7908 11336 7936
rect 11330 7896 11336 7908
rect 11388 7936 11394 7948
rect 12268 7936 12296 8032
rect 11388 7908 12296 7936
rect 11388 7896 11394 7908
rect 16574 7896 16580 7948
rect 16632 7936 16638 7948
rect 17221 7939 17279 7945
rect 17221 7936 17233 7939
rect 16632 7908 17233 7936
rect 16632 7896 16638 7908
rect 17221 7905 17233 7908
rect 17267 7905 17279 7939
rect 17221 7899 17279 7905
rect 9493 7871 9551 7877
rect 9493 7837 9505 7871
rect 9539 7868 9551 7871
rect 10318 7868 10324 7880
rect 9539 7840 10324 7868
rect 9539 7837 9551 7840
rect 9493 7831 9551 7837
rect 10318 7828 10324 7840
rect 10376 7828 10382 7880
rect 11514 7868 11520 7880
rect 11475 7840 11520 7868
rect 11514 7828 11520 7840
rect 11572 7828 11578 7880
rect 12345 7871 12403 7877
rect 12345 7837 12357 7871
rect 12391 7868 12403 7871
rect 12526 7868 12532 7880
rect 12391 7840 12532 7868
rect 12391 7837 12403 7840
rect 12345 7831 12403 7837
rect 12526 7828 12532 7840
rect 12584 7828 12590 7880
rect 17310 7828 17316 7880
rect 17368 7868 17374 7880
rect 17477 7871 17535 7877
rect 17477 7868 17489 7871
rect 17368 7840 17489 7868
rect 17368 7828 17374 7840
rect 17477 7837 17489 7840
rect 17523 7837 17535 7871
rect 17477 7831 17535 7837
rect 9766 7809 9772 7812
rect 9760 7763 9772 7809
rect 9824 7800 9830 7812
rect 9824 7772 9860 7800
rect 9766 7760 9772 7763
rect 9824 7760 9830 7772
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 9766 7528 9772 7540
rect 9727 7500 9772 7528
rect 9766 7488 9772 7500
rect 9824 7488 9830 7540
rect 17586 7528 17592 7540
rect 17547 7500 17592 7528
rect 17586 7488 17592 7500
rect 17644 7488 17650 7540
rect 9950 7392 9956 7404
rect 9911 7364 9956 7392
rect 9950 7352 9956 7364
rect 10008 7352 10014 7404
rect 17218 7392 17224 7404
rect 17179 7364 17224 7392
rect 17218 7352 17224 7364
rect 17276 7352 17282 7404
rect 17402 7392 17408 7404
rect 17363 7364 17408 7392
rect 17402 7352 17408 7364
rect 17460 7352 17466 7404
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 9033 6851 9091 6857
rect 9033 6817 9045 6851
rect 9079 6848 9091 6851
rect 9401 6851 9459 6857
rect 9079 6820 9352 6848
rect 9079 6817 9091 6820
rect 9033 6811 9091 6817
rect 9214 6780 9220 6792
rect 9175 6752 9220 6780
rect 9214 6740 9220 6752
rect 9272 6740 9278 6792
rect 9324 6780 9352 6820
rect 9401 6817 9413 6851
rect 9447 6848 9459 6851
rect 9950 6848 9956 6860
rect 9447 6820 9956 6848
rect 9447 6817 9459 6820
rect 9401 6811 9459 6817
rect 9950 6808 9956 6820
rect 10008 6808 10014 6860
rect 11330 6780 11336 6792
rect 9324 6752 11336 6780
rect 11330 6740 11336 6752
rect 11388 6740 11394 6792
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 1397 2635 1455 2641
rect 1397 2601 1409 2635
rect 1443 2632 1455 2635
rect 9214 2632 9220 2644
rect 1443 2604 9220 2632
rect 1443 2601 1455 2604
rect 1397 2595 1455 2601
rect 9214 2592 9220 2604
rect 9272 2592 9278 2644
rect 10413 2635 10471 2641
rect 10413 2601 10425 2635
rect 10459 2632 10471 2635
rect 11238 2632 11244 2644
rect 10459 2604 11244 2632
rect 10459 2601 10471 2604
rect 10413 2595 10471 2601
rect 11238 2592 11244 2604
rect 11296 2592 11302 2644
rect 17402 2456 17408 2508
rect 17460 2496 17466 2508
rect 31021 2499 31079 2505
rect 31021 2496 31033 2499
rect 17460 2468 31033 2496
rect 17460 2456 17466 2468
rect 31021 2465 31033 2468
rect 31067 2465 31079 2499
rect 31021 2459 31079 2465
rect 14 2388 20 2440
rect 72 2428 78 2440
rect 1581 2431 1639 2437
rect 1581 2428 1593 2431
rect 72 2400 1593 2428
rect 72 2388 78 2400
rect 1581 2397 1593 2400
rect 1627 2397 1639 2431
rect 1581 2391 1639 2397
rect 10318 2388 10324 2440
rect 10376 2428 10382 2440
rect 10597 2431 10655 2437
rect 10597 2428 10609 2431
rect 10376 2400 10609 2428
rect 10376 2388 10382 2400
rect 10597 2397 10609 2400
rect 10643 2397 10655 2431
rect 10597 2391 10655 2397
rect 20717 2431 20775 2437
rect 20717 2397 20729 2431
rect 20763 2428 20775 2431
rect 26510 2428 26516 2440
rect 20763 2400 26516 2428
rect 20763 2397 20775 2400
rect 20717 2391 20775 2397
rect 26510 2388 26516 2400
rect 26568 2388 26574 2440
rect 30745 2431 30803 2437
rect 30745 2397 30757 2431
rect 30791 2428 30803 2431
rect 30926 2428 30932 2440
rect 30791 2400 30932 2428
rect 30791 2397 30803 2400
rect 30745 2391 30803 2397
rect 30926 2388 30932 2400
rect 30984 2388 30990 2440
rect 37734 2388 37740 2440
rect 37792 2428 37798 2440
rect 37829 2431 37887 2437
rect 37829 2428 37841 2431
rect 37792 2400 37841 2428
rect 37792 2388 37798 2400
rect 37829 2397 37841 2400
rect 37875 2397 37887 2431
rect 37829 2391 37887 2397
rect 20622 2252 20628 2304
rect 20680 2292 20686 2304
rect 20901 2295 20959 2301
rect 20901 2292 20913 2295
rect 20680 2264 20913 2292
rect 20680 2252 20686 2264
rect 20901 2261 20913 2264
rect 20947 2261 20959 2295
rect 38010 2292 38016 2304
rect 37971 2264 38016 2292
rect 20901 2255 20959 2261
rect 38010 2252 38016 2264
rect 38068 2252 38074 2304
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 25228 37451 25280 37460
rect 25228 37417 25237 37451
rect 25237 37417 25271 37451
rect 25271 37417 25280 37451
rect 25228 37408 25280 37417
rect 24492 37340 24544 37392
rect 25504 37340 25556 37392
rect 25872 37383 25924 37392
rect 25872 37349 25881 37383
rect 25881 37349 25915 37383
rect 25915 37349 25924 37383
rect 25872 37340 25924 37349
rect 3792 37247 3844 37256
rect 3792 37213 3801 37247
rect 3801 37213 3835 37247
rect 3835 37213 3844 37247
rect 3792 37204 3844 37213
rect 14924 37204 14976 37256
rect 23848 37204 23900 37256
rect 25412 37247 25464 37256
rect 25412 37213 25421 37247
rect 25421 37213 25455 37247
rect 25455 37213 25464 37247
rect 27620 37272 27672 37324
rect 25412 37204 25464 37213
rect 26424 37204 26476 37256
rect 28632 37247 28684 37256
rect 26976 37179 27028 37188
rect 26976 37145 26985 37179
rect 26985 37145 27019 37179
rect 27019 37145 27028 37179
rect 26976 37136 27028 37145
rect 28264 37179 28316 37188
rect 3240 37068 3292 37120
rect 13544 37068 13596 37120
rect 26332 37068 26384 37120
rect 26424 37068 26476 37120
rect 28264 37145 28273 37179
rect 28273 37145 28307 37179
rect 28307 37145 28316 37179
rect 28264 37136 28316 37145
rect 28632 37213 28641 37247
rect 28641 37213 28675 37247
rect 28675 37213 28684 37247
rect 30288 37247 30340 37256
rect 28632 37204 28684 37213
rect 30288 37213 30297 37247
rect 30297 37213 30331 37247
rect 30331 37213 30340 37247
rect 30288 37204 30340 37213
rect 29736 37136 29788 37188
rect 35808 37204 35860 37256
rect 28816 37068 28868 37120
rect 30472 37068 30524 37120
rect 34520 37068 34572 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 25228 36864 25280 36916
rect 28816 36907 28868 36916
rect 28816 36873 28825 36907
rect 28825 36873 28859 36907
rect 28859 36873 28868 36907
rect 28816 36864 28868 36873
rect 29644 36864 29696 36916
rect 24400 36839 24452 36848
rect 24400 36805 24409 36839
rect 24409 36805 24443 36839
rect 24443 36805 24452 36839
rect 24400 36796 24452 36805
rect 28264 36796 28316 36848
rect 24308 36728 24360 36780
rect 24768 36728 24820 36780
rect 25504 36592 25556 36644
rect 24952 36567 25004 36576
rect 24952 36533 24961 36567
rect 24961 36533 24995 36567
rect 24995 36533 25004 36567
rect 24952 36524 25004 36533
rect 26240 36660 26292 36712
rect 27620 36728 27672 36780
rect 28632 36771 28684 36780
rect 28632 36737 28641 36771
rect 28641 36737 28675 36771
rect 28675 36737 28684 36771
rect 28632 36728 28684 36737
rect 29736 36728 29788 36780
rect 29828 36771 29880 36780
rect 29828 36737 29837 36771
rect 29837 36737 29871 36771
rect 29871 36737 29880 36771
rect 30472 36771 30524 36780
rect 29828 36728 29880 36737
rect 30472 36737 30481 36771
rect 30481 36737 30515 36771
rect 30515 36737 30524 36771
rect 30472 36728 30524 36737
rect 30196 36660 30248 36712
rect 26332 36592 26384 36644
rect 30380 36592 30432 36644
rect 30932 36660 30984 36712
rect 32496 36592 32548 36644
rect 27528 36524 27580 36576
rect 27712 36567 27764 36576
rect 27712 36533 27721 36567
rect 27721 36533 27755 36567
rect 27755 36533 27764 36567
rect 27712 36524 27764 36533
rect 28908 36524 28960 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 24400 36320 24452 36372
rect 26056 36320 26108 36372
rect 26240 36363 26292 36372
rect 26240 36329 26249 36363
rect 26249 36329 26283 36363
rect 26283 36329 26292 36363
rect 26240 36320 26292 36329
rect 26976 36320 27028 36372
rect 27528 36320 27580 36372
rect 28816 36320 28868 36372
rect 25412 36252 25464 36304
rect 28908 36252 28960 36304
rect 30932 36363 30984 36372
rect 28816 36227 28868 36236
rect 28816 36193 28825 36227
rect 28825 36193 28859 36227
rect 28859 36193 28868 36227
rect 30288 36252 30340 36304
rect 30932 36329 30941 36363
rect 30941 36329 30975 36363
rect 30975 36329 30984 36363
rect 30932 36320 30984 36329
rect 31576 36363 31628 36372
rect 31576 36329 31585 36363
rect 31585 36329 31619 36363
rect 31619 36329 31628 36363
rect 31576 36320 31628 36329
rect 28816 36184 28868 36193
rect 25044 36116 25096 36168
rect 25872 36116 25924 36168
rect 26424 36159 26476 36168
rect 26424 36125 26433 36159
rect 26433 36125 26467 36159
rect 26467 36125 26476 36159
rect 26424 36116 26476 36125
rect 29644 36159 29696 36168
rect 29644 36125 29653 36159
rect 29653 36125 29687 36159
rect 29687 36125 29696 36159
rect 29644 36116 29696 36125
rect 24308 36048 24360 36100
rect 30196 36116 30248 36168
rect 31208 36116 31260 36168
rect 24860 35980 24912 36032
rect 31300 36048 31352 36100
rect 32128 36184 32180 36236
rect 31668 36159 31720 36168
rect 31668 36125 31677 36159
rect 31677 36125 31711 36159
rect 31711 36125 31720 36159
rect 31668 36116 31720 36125
rect 32220 36116 32272 36168
rect 32404 36159 32456 36168
rect 32404 36125 32413 36159
rect 32413 36125 32447 36159
rect 32447 36125 32456 36159
rect 32404 36116 32456 36125
rect 28264 36023 28316 36032
rect 28264 35989 28273 36023
rect 28273 35989 28307 36023
rect 28307 35989 28316 36023
rect 28264 35980 28316 35989
rect 28632 36023 28684 36032
rect 28632 35989 28641 36023
rect 28641 35989 28675 36023
rect 28675 35989 28684 36023
rect 28632 35980 28684 35989
rect 30288 35980 30340 36032
rect 31852 36023 31904 36032
rect 31852 35989 31861 36023
rect 31861 35989 31895 36023
rect 31895 35989 31904 36023
rect 31852 35980 31904 35989
rect 32956 35980 33008 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 24768 35819 24820 35828
rect 24768 35785 24777 35819
rect 24777 35785 24811 35819
rect 24811 35785 24820 35819
rect 24768 35776 24820 35785
rect 26148 35776 26200 35828
rect 27712 35776 27764 35828
rect 23756 35683 23808 35692
rect 23756 35649 23765 35683
rect 23765 35649 23799 35683
rect 23799 35649 23808 35683
rect 23756 35640 23808 35649
rect 24400 35640 24452 35692
rect 24032 35572 24084 35624
rect 25320 35683 25372 35692
rect 25320 35649 25329 35683
rect 25329 35649 25363 35683
rect 25363 35649 25372 35683
rect 25320 35640 25372 35649
rect 25412 35572 25464 35624
rect 28540 35776 28592 35828
rect 29736 35776 29788 35828
rect 30288 35776 30340 35828
rect 32496 35819 32548 35828
rect 32496 35785 32505 35819
rect 32505 35785 32539 35819
rect 32539 35785 32548 35819
rect 32496 35776 32548 35785
rect 28724 35751 28776 35760
rect 26332 35640 26384 35692
rect 26792 35640 26844 35692
rect 28724 35717 28733 35751
rect 28733 35717 28767 35751
rect 28767 35717 28776 35751
rect 28724 35708 28776 35717
rect 28448 35683 28500 35692
rect 28448 35649 28457 35683
rect 28457 35649 28491 35683
rect 28491 35649 28500 35683
rect 28448 35640 28500 35649
rect 26516 35572 26568 35624
rect 27528 35615 27580 35624
rect 27528 35581 27537 35615
rect 27537 35581 27571 35615
rect 27571 35581 27580 35615
rect 27528 35572 27580 35581
rect 28356 35572 28408 35624
rect 30380 35640 30432 35692
rect 31300 35683 31352 35692
rect 31300 35649 31309 35683
rect 31309 35649 31343 35683
rect 31343 35649 31352 35683
rect 31300 35640 31352 35649
rect 32128 35683 32180 35692
rect 31852 35572 31904 35624
rect 32128 35649 32137 35683
rect 32137 35649 32171 35683
rect 32171 35649 32180 35683
rect 32128 35640 32180 35649
rect 32956 35683 33008 35692
rect 32956 35649 32965 35683
rect 32965 35649 32999 35683
rect 32999 35649 33008 35683
rect 32956 35640 33008 35649
rect 32220 35615 32272 35624
rect 32220 35581 32229 35615
rect 32229 35581 32263 35615
rect 32263 35581 32272 35615
rect 32220 35572 32272 35581
rect 23848 35504 23900 35556
rect 28172 35504 28224 35556
rect 23664 35479 23716 35488
rect 23664 35445 23673 35479
rect 23673 35445 23707 35479
rect 23707 35445 23716 35479
rect 23664 35436 23716 35445
rect 27252 35436 27304 35488
rect 28448 35436 28500 35488
rect 31300 35436 31352 35488
rect 32496 35436 32548 35488
rect 33048 35479 33100 35488
rect 33048 35445 33057 35479
rect 33057 35445 33091 35479
rect 33091 35445 33100 35479
rect 33048 35436 33100 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 24400 35275 24452 35284
rect 24400 35241 24409 35275
rect 24409 35241 24443 35275
rect 24443 35241 24452 35275
rect 24400 35232 24452 35241
rect 25320 35232 25372 35284
rect 28632 35275 28684 35284
rect 28632 35241 28641 35275
rect 28641 35241 28675 35275
rect 28675 35241 28684 35275
rect 28632 35232 28684 35241
rect 29828 35232 29880 35284
rect 31668 35232 31720 35284
rect 32128 35232 32180 35284
rect 26424 35164 26476 35216
rect 27804 35207 27856 35216
rect 27804 35173 27813 35207
rect 27813 35173 27847 35207
rect 27847 35173 27856 35207
rect 27804 35164 27856 35173
rect 20168 35071 20220 35080
rect 20168 35037 20177 35071
rect 20177 35037 20211 35071
rect 20211 35037 20220 35071
rect 20168 35028 20220 35037
rect 20444 35028 20496 35080
rect 20812 35071 20864 35080
rect 20812 35037 20821 35071
rect 20821 35037 20855 35071
rect 20855 35037 20864 35071
rect 20812 35028 20864 35037
rect 20996 35071 21048 35080
rect 20996 35037 21005 35071
rect 21005 35037 21039 35071
rect 21039 35037 21048 35071
rect 20996 35028 21048 35037
rect 21824 35028 21876 35080
rect 27620 35096 27672 35148
rect 28816 35096 28868 35148
rect 30932 35139 30984 35148
rect 30932 35105 30941 35139
rect 30941 35105 30975 35139
rect 30975 35105 30984 35139
rect 30932 35096 30984 35105
rect 33048 35164 33100 35216
rect 23848 35071 23900 35080
rect 23848 35037 23857 35071
rect 23857 35037 23891 35071
rect 23891 35037 23900 35071
rect 23848 35028 23900 35037
rect 24032 35028 24084 35080
rect 24400 35028 24452 35080
rect 23756 34960 23808 35012
rect 25504 35028 25556 35080
rect 25688 35028 25740 35080
rect 26148 35028 26200 35080
rect 26424 35028 26476 35080
rect 26608 35028 26660 35080
rect 27896 35028 27948 35080
rect 28080 35071 28132 35080
rect 28080 35037 28089 35071
rect 28089 35037 28123 35071
rect 28123 35037 28132 35071
rect 28080 35028 28132 35037
rect 28540 35071 28592 35080
rect 28540 35037 28549 35071
rect 28549 35037 28583 35071
rect 28583 35037 28592 35071
rect 28540 35028 28592 35037
rect 26332 34960 26384 35012
rect 26976 34960 27028 35012
rect 20260 34935 20312 34944
rect 20260 34901 20269 34935
rect 20269 34901 20303 34935
rect 20303 34901 20312 34935
rect 20260 34892 20312 34901
rect 20352 34892 20404 34944
rect 24676 34892 24728 34944
rect 24768 34892 24820 34944
rect 26424 34892 26476 34944
rect 26792 34892 26844 34944
rect 28448 34960 28500 35012
rect 30288 35028 30340 35080
rect 30380 35028 30432 35080
rect 31576 35071 31628 35080
rect 31576 35037 31585 35071
rect 31585 35037 31619 35071
rect 31619 35037 31628 35071
rect 31576 35028 31628 35037
rect 31668 35028 31720 35080
rect 27988 34935 28040 34944
rect 27988 34901 27997 34935
rect 27997 34901 28031 34935
rect 28031 34901 28040 34935
rect 27988 34892 28040 34901
rect 28172 34892 28224 34944
rect 29736 34892 29788 34944
rect 30196 34892 30248 34944
rect 30472 34892 30524 34944
rect 31392 34892 31444 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 20812 34688 20864 34740
rect 21824 34731 21876 34740
rect 21824 34697 21833 34731
rect 21833 34697 21867 34731
rect 21867 34697 21876 34731
rect 21824 34688 21876 34697
rect 26148 34688 26200 34740
rect 26424 34620 26476 34672
rect 19984 34552 20036 34604
rect 20260 34595 20312 34604
rect 20260 34561 20269 34595
rect 20269 34561 20303 34595
rect 20303 34561 20312 34595
rect 20260 34552 20312 34561
rect 21088 34595 21140 34604
rect 21088 34561 21097 34595
rect 21097 34561 21131 34595
rect 21131 34561 21140 34595
rect 21088 34552 21140 34561
rect 23664 34552 23716 34604
rect 24676 34552 24728 34604
rect 24860 34595 24912 34604
rect 24860 34561 24869 34595
rect 24869 34561 24903 34595
rect 24903 34561 24912 34595
rect 24860 34552 24912 34561
rect 25320 34552 25372 34604
rect 25872 34552 25924 34604
rect 26516 34552 26568 34604
rect 20352 34527 20404 34536
rect 20352 34493 20361 34527
rect 20361 34493 20395 34527
rect 20395 34493 20404 34527
rect 20352 34484 20404 34493
rect 23572 34527 23624 34536
rect 23572 34493 23581 34527
rect 23581 34493 23615 34527
rect 23615 34493 23624 34527
rect 23572 34484 23624 34493
rect 23756 34484 23808 34536
rect 26884 34552 26936 34604
rect 27712 34620 27764 34672
rect 27896 34688 27948 34740
rect 31392 34731 31444 34740
rect 27988 34620 28040 34672
rect 28540 34620 28592 34672
rect 30196 34663 30248 34672
rect 30196 34629 30205 34663
rect 30205 34629 30239 34663
rect 30239 34629 30248 34663
rect 30196 34620 30248 34629
rect 30288 34620 30340 34672
rect 31392 34697 31401 34731
rect 31401 34697 31435 34731
rect 31435 34697 31444 34731
rect 31392 34688 31444 34697
rect 27620 34595 27672 34604
rect 27620 34561 27629 34595
rect 27629 34561 27663 34595
rect 27663 34561 27672 34595
rect 27620 34552 27672 34561
rect 28172 34552 28224 34604
rect 29276 34595 29328 34604
rect 29276 34561 29285 34595
rect 29285 34561 29319 34595
rect 29319 34561 29328 34595
rect 29276 34552 29328 34561
rect 29460 34595 29512 34604
rect 29460 34561 29469 34595
rect 29469 34561 29503 34595
rect 29503 34561 29512 34595
rect 29460 34552 29512 34561
rect 31024 34595 31076 34604
rect 31024 34561 31033 34595
rect 31033 34561 31067 34595
rect 31067 34561 31076 34595
rect 31024 34552 31076 34561
rect 31576 34620 31628 34672
rect 34612 34620 34664 34672
rect 32220 34552 32272 34604
rect 38200 34552 38252 34604
rect 32404 34527 32456 34536
rect 32404 34493 32413 34527
rect 32413 34493 32447 34527
rect 32447 34493 32456 34527
rect 32404 34484 32456 34493
rect 22836 34416 22888 34468
rect 24032 34416 24084 34468
rect 28080 34348 28132 34400
rect 28632 34391 28684 34400
rect 28632 34357 28641 34391
rect 28641 34357 28675 34391
rect 28675 34357 28684 34391
rect 28632 34348 28684 34357
rect 28816 34391 28868 34400
rect 28816 34357 28825 34391
rect 28825 34357 28859 34391
rect 28859 34357 28868 34391
rect 28816 34348 28868 34357
rect 29828 34348 29880 34400
rect 30380 34391 30432 34400
rect 30380 34357 30389 34391
rect 30389 34357 30423 34391
rect 30423 34357 30432 34391
rect 30380 34348 30432 34357
rect 31024 34348 31076 34400
rect 31392 34348 31444 34400
rect 31760 34348 31812 34400
rect 32312 34391 32364 34400
rect 32312 34357 32321 34391
rect 32321 34357 32355 34391
rect 32355 34357 32364 34391
rect 38016 34391 38068 34400
rect 32312 34348 32364 34357
rect 38016 34357 38025 34391
rect 38025 34357 38059 34391
rect 38059 34357 38068 34391
rect 38016 34348 38068 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 21088 34144 21140 34196
rect 25596 34144 25648 34196
rect 20076 34076 20128 34128
rect 20996 34008 21048 34060
rect 19248 33940 19300 33992
rect 19984 33940 20036 33992
rect 20260 33940 20312 33992
rect 20812 33983 20864 33992
rect 20812 33949 20821 33983
rect 20821 33949 20855 33983
rect 20855 33949 20864 33983
rect 20812 33940 20864 33949
rect 28448 34144 28500 34196
rect 29644 34144 29696 34196
rect 29920 34144 29972 34196
rect 30288 34144 30340 34196
rect 31392 34144 31444 34196
rect 23572 34008 23624 34060
rect 24124 34008 24176 34060
rect 24768 34008 24820 34060
rect 25504 34051 25556 34060
rect 23480 33983 23532 33992
rect 23480 33949 23489 33983
rect 23489 33949 23523 33983
rect 23523 33949 23532 33983
rect 23480 33940 23532 33949
rect 23756 33983 23808 33992
rect 23756 33949 23765 33983
rect 23765 33949 23799 33983
rect 23799 33949 23808 33983
rect 23756 33940 23808 33949
rect 24860 33983 24912 33992
rect 23940 33872 23992 33924
rect 24400 33872 24452 33924
rect 24860 33949 24869 33983
rect 24869 33949 24903 33983
rect 24903 33949 24912 33983
rect 24860 33940 24912 33949
rect 25504 34017 25513 34051
rect 25513 34017 25547 34051
rect 25547 34017 25556 34051
rect 25504 34008 25556 34017
rect 25964 33983 26016 33992
rect 25964 33949 25973 33983
rect 25973 33949 26007 33983
rect 26007 33949 26016 33983
rect 25964 33940 26016 33949
rect 26516 33940 26568 33992
rect 27436 33940 27488 33992
rect 27804 33940 27856 33992
rect 28816 34008 28868 34060
rect 31668 34076 31720 34128
rect 31944 34076 31996 34128
rect 29644 34051 29696 34060
rect 29644 34017 29653 34051
rect 29653 34017 29687 34051
rect 29687 34017 29696 34051
rect 29644 34008 29696 34017
rect 29828 33983 29880 33992
rect 29828 33949 29837 33983
rect 29837 33949 29871 33983
rect 29871 33949 29880 33983
rect 29828 33940 29880 33949
rect 28724 33872 28776 33924
rect 30288 33872 30340 33924
rect 30748 33940 30800 33992
rect 32404 34008 32456 34060
rect 33048 34051 33100 34060
rect 33048 34017 33057 34051
rect 33057 34017 33091 34051
rect 33091 34017 33100 34051
rect 33048 34008 33100 34017
rect 31944 33983 31996 33992
rect 31944 33949 31953 33983
rect 31953 33949 31987 33983
rect 31987 33949 31996 33983
rect 31944 33940 31996 33949
rect 32772 33983 32824 33992
rect 20352 33804 20404 33856
rect 20720 33847 20772 33856
rect 20720 33813 20729 33847
rect 20729 33813 20763 33847
rect 20763 33813 20772 33847
rect 20720 33804 20772 33813
rect 30196 33804 30248 33856
rect 30840 33804 30892 33856
rect 31208 33804 31260 33856
rect 32220 33872 32272 33924
rect 32772 33949 32781 33983
rect 32781 33949 32815 33983
rect 32815 33949 32824 33983
rect 32772 33940 32824 33949
rect 33876 33940 33928 33992
rect 32680 33872 32732 33924
rect 31668 33804 31720 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 20996 33600 21048 33652
rect 19432 33464 19484 33516
rect 20076 33464 20128 33516
rect 20260 33507 20312 33516
rect 20260 33473 20269 33507
rect 20269 33473 20303 33507
rect 20303 33473 20312 33507
rect 20260 33464 20312 33473
rect 20352 33507 20404 33516
rect 20352 33473 20361 33507
rect 20361 33473 20395 33507
rect 20395 33473 20404 33507
rect 20812 33532 20864 33584
rect 24124 33575 24176 33584
rect 24124 33541 24133 33575
rect 24133 33541 24167 33575
rect 24167 33541 24176 33575
rect 24124 33532 24176 33541
rect 25964 33600 26016 33652
rect 26976 33643 27028 33652
rect 26976 33609 26985 33643
rect 26985 33609 27019 33643
rect 27019 33609 27028 33643
rect 26976 33600 27028 33609
rect 30288 33643 30340 33652
rect 30288 33609 30297 33643
rect 30297 33609 30331 33643
rect 30331 33609 30340 33643
rect 30288 33600 30340 33609
rect 20352 33464 20404 33473
rect 22192 33507 22244 33516
rect 19984 33396 20036 33448
rect 20444 33396 20496 33448
rect 22192 33473 22201 33507
rect 22201 33473 22235 33507
rect 22235 33473 22244 33507
rect 22192 33464 22244 33473
rect 23940 33507 23992 33516
rect 23940 33473 23949 33507
rect 23949 33473 23983 33507
rect 23983 33473 23992 33507
rect 23940 33464 23992 33473
rect 24032 33507 24084 33516
rect 24032 33473 24041 33507
rect 24041 33473 24075 33507
rect 24075 33473 24084 33507
rect 29276 33532 29328 33584
rect 31208 33575 31260 33584
rect 24032 33464 24084 33473
rect 24860 33507 24912 33516
rect 20812 33396 20864 33448
rect 22284 33439 22336 33448
rect 22284 33405 22293 33439
rect 22293 33405 22327 33439
rect 22327 33405 22336 33439
rect 22284 33396 22336 33405
rect 22836 33396 22888 33448
rect 23480 33396 23532 33448
rect 24860 33473 24869 33507
rect 24869 33473 24903 33507
rect 24903 33473 24912 33507
rect 24860 33464 24912 33473
rect 25780 33464 25832 33516
rect 25872 33507 25924 33516
rect 25872 33473 25881 33507
rect 25881 33473 25915 33507
rect 25915 33473 25924 33507
rect 25872 33464 25924 33473
rect 26056 33464 26108 33516
rect 27436 33507 27488 33516
rect 27436 33473 27445 33507
rect 27445 33473 27479 33507
rect 27479 33473 27488 33507
rect 27436 33464 27488 33473
rect 28448 33507 28500 33516
rect 28448 33473 28457 33507
rect 28457 33473 28491 33507
rect 28491 33473 28500 33507
rect 28448 33464 28500 33473
rect 28632 33464 28684 33516
rect 29092 33507 29144 33516
rect 29092 33473 29101 33507
rect 29101 33473 29135 33507
rect 29135 33473 29144 33507
rect 29092 33464 29144 33473
rect 29460 33464 29512 33516
rect 31208 33541 31217 33575
rect 31217 33541 31251 33575
rect 31251 33541 31260 33575
rect 31208 33532 31260 33541
rect 31668 33532 31720 33584
rect 32772 33532 32824 33584
rect 31300 33507 31352 33516
rect 24676 33396 24728 33448
rect 25504 33396 25556 33448
rect 25596 33439 25648 33448
rect 25596 33405 25605 33439
rect 25605 33405 25639 33439
rect 25639 33405 25648 33439
rect 25596 33396 25648 33405
rect 29000 33396 29052 33448
rect 24860 33328 24912 33380
rect 25044 33328 25096 33380
rect 28724 33371 28776 33380
rect 28724 33337 28733 33371
rect 28733 33337 28767 33371
rect 28767 33337 28776 33371
rect 28724 33328 28776 33337
rect 31300 33473 31309 33507
rect 31309 33473 31343 33507
rect 31343 33473 31352 33507
rect 31300 33464 31352 33473
rect 31392 33507 31444 33516
rect 31392 33473 31425 33507
rect 31425 33473 31444 33507
rect 31392 33464 31444 33473
rect 31944 33464 31996 33516
rect 32864 33464 32916 33516
rect 32312 33396 32364 33448
rect 33876 33439 33928 33448
rect 18328 33260 18380 33312
rect 19248 33260 19300 33312
rect 21088 33260 21140 33312
rect 23664 33260 23716 33312
rect 24400 33260 24452 33312
rect 31300 33260 31352 33312
rect 31852 33328 31904 33380
rect 33876 33405 33885 33439
rect 33885 33405 33919 33439
rect 33919 33405 33928 33439
rect 33876 33396 33928 33405
rect 34796 33328 34848 33380
rect 32588 33260 32640 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 20812 33056 20864 33108
rect 23756 33056 23808 33108
rect 25596 33056 25648 33108
rect 26240 33056 26292 33108
rect 28540 33056 28592 33108
rect 1492 32852 1544 32904
rect 16764 32895 16816 32904
rect 16764 32861 16773 32895
rect 16773 32861 16807 32895
rect 16807 32861 16816 32895
rect 16764 32852 16816 32861
rect 16856 32852 16908 32904
rect 17224 32895 17276 32904
rect 17224 32861 17233 32895
rect 17233 32861 17267 32895
rect 17267 32861 17276 32895
rect 17224 32852 17276 32861
rect 18052 32895 18104 32904
rect 18052 32861 18061 32895
rect 18061 32861 18095 32895
rect 18095 32861 18104 32895
rect 18052 32852 18104 32861
rect 20720 32852 20772 32904
rect 22284 32988 22336 33040
rect 24676 33031 24728 33040
rect 24676 32997 24685 33031
rect 24685 32997 24719 33031
rect 24719 32997 24728 33031
rect 24676 32988 24728 32997
rect 23756 32920 23808 32972
rect 22192 32852 22244 32904
rect 23664 32895 23716 32904
rect 23664 32861 23673 32895
rect 23673 32861 23707 32895
rect 23707 32861 23716 32895
rect 23664 32852 23716 32861
rect 24676 32895 24728 32904
rect 24676 32861 24685 32895
rect 24685 32861 24719 32895
rect 24719 32861 24728 32895
rect 24676 32852 24728 32861
rect 25228 32895 25280 32904
rect 25228 32861 25237 32895
rect 25237 32861 25271 32895
rect 25271 32861 25280 32895
rect 25228 32852 25280 32861
rect 26516 32988 26568 33040
rect 25872 32920 25924 32972
rect 26424 32920 26476 32972
rect 1584 32759 1636 32768
rect 1584 32725 1593 32759
rect 1593 32725 1627 32759
rect 1627 32725 1636 32759
rect 1584 32716 1636 32725
rect 17316 32716 17368 32768
rect 24124 32784 24176 32836
rect 24860 32784 24912 32836
rect 26332 32895 26384 32904
rect 26332 32861 26341 32895
rect 26341 32861 26375 32895
rect 26375 32861 26384 32895
rect 26332 32852 26384 32861
rect 25780 32784 25832 32836
rect 18144 32759 18196 32768
rect 18144 32725 18153 32759
rect 18153 32725 18187 32759
rect 18187 32725 18196 32759
rect 18144 32716 18196 32725
rect 21916 32716 21968 32768
rect 23204 32716 23256 32768
rect 27436 32895 27488 32904
rect 27436 32861 27445 32895
rect 27445 32861 27479 32895
rect 27479 32861 27488 32895
rect 27436 32852 27488 32861
rect 29092 32920 29144 32972
rect 29644 32920 29696 32972
rect 31208 32988 31260 33040
rect 30380 32920 30432 32972
rect 30932 32920 30984 32972
rect 32496 33056 32548 33108
rect 31760 32988 31812 33040
rect 33416 32988 33468 33040
rect 27344 32759 27396 32768
rect 27344 32725 27353 32759
rect 27353 32725 27387 32759
rect 27387 32725 27396 32759
rect 27344 32716 27396 32725
rect 27620 32784 27672 32836
rect 28448 32784 28500 32836
rect 29000 32852 29052 32904
rect 29920 32852 29972 32904
rect 31852 32895 31904 32904
rect 30656 32784 30708 32836
rect 31484 32784 31536 32836
rect 31852 32861 31861 32895
rect 31861 32861 31895 32895
rect 31895 32861 31904 32895
rect 31852 32852 31904 32861
rect 33048 32920 33100 32972
rect 34796 32963 34848 32972
rect 34796 32929 34805 32963
rect 34805 32929 34839 32963
rect 34839 32929 34848 32963
rect 34796 32920 34848 32929
rect 32496 32895 32548 32904
rect 32496 32861 32505 32895
rect 32505 32861 32539 32895
rect 32539 32861 32548 32895
rect 32496 32852 32548 32861
rect 31760 32784 31812 32836
rect 31944 32784 31996 32836
rect 32680 32895 32732 32904
rect 32680 32861 32689 32895
rect 32689 32861 32723 32895
rect 32723 32861 32732 32895
rect 32864 32895 32916 32904
rect 32680 32852 32732 32861
rect 32864 32861 32873 32895
rect 32873 32861 32907 32895
rect 32907 32861 32916 32895
rect 32864 32852 32916 32861
rect 32956 32852 33008 32904
rect 32772 32784 32824 32836
rect 33968 32895 34020 32904
rect 33968 32861 33977 32895
rect 33977 32861 34011 32895
rect 34011 32861 34020 32895
rect 33968 32852 34020 32861
rect 28172 32716 28224 32768
rect 28540 32716 28592 32768
rect 30748 32716 30800 32768
rect 33784 32716 33836 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 16304 32376 16356 32428
rect 16764 32376 16816 32428
rect 17316 32419 17368 32428
rect 17316 32385 17325 32419
rect 17325 32385 17359 32419
rect 17359 32385 17368 32419
rect 17316 32376 17368 32385
rect 15292 32308 15344 32360
rect 17224 32351 17276 32360
rect 17224 32317 17233 32351
rect 17233 32317 17267 32351
rect 17267 32317 17276 32351
rect 17224 32308 17276 32317
rect 19064 32512 19116 32564
rect 21088 32555 21140 32564
rect 21088 32521 21113 32555
rect 21113 32521 21140 32555
rect 21088 32512 21140 32521
rect 18144 32376 18196 32428
rect 20812 32444 20864 32496
rect 22284 32444 22336 32496
rect 23664 32512 23716 32564
rect 24676 32512 24728 32564
rect 18972 32376 19024 32428
rect 19156 32376 19208 32428
rect 19984 32308 20036 32360
rect 16856 32240 16908 32292
rect 19248 32240 19300 32292
rect 22836 32419 22888 32428
rect 22836 32385 22845 32419
rect 22845 32385 22879 32419
rect 22879 32385 22888 32419
rect 22836 32376 22888 32385
rect 23020 32419 23072 32428
rect 23020 32385 23029 32419
rect 23029 32385 23063 32419
rect 23063 32385 23072 32419
rect 23020 32376 23072 32385
rect 23572 32376 23624 32428
rect 25228 32444 25280 32496
rect 23756 32308 23808 32360
rect 24860 32308 24912 32360
rect 25780 32376 25832 32428
rect 26332 32512 26384 32564
rect 27160 32512 27212 32564
rect 28540 32512 28592 32564
rect 29000 32512 29052 32564
rect 27344 32487 27396 32496
rect 26056 32376 26108 32428
rect 27344 32453 27353 32487
rect 27353 32453 27387 32487
rect 27387 32453 27396 32487
rect 27344 32444 27396 32453
rect 31576 32512 31628 32564
rect 31668 32512 31720 32564
rect 30472 32487 30524 32496
rect 30472 32453 30507 32487
rect 30507 32453 30524 32487
rect 30472 32444 30524 32453
rect 31392 32444 31444 32496
rect 25044 32240 25096 32292
rect 26700 32376 26752 32428
rect 27160 32419 27212 32428
rect 27160 32385 27169 32419
rect 27169 32385 27203 32419
rect 27203 32385 27212 32419
rect 27160 32376 27212 32385
rect 27436 32419 27488 32428
rect 27436 32385 27445 32419
rect 27445 32385 27479 32419
rect 27479 32385 27488 32419
rect 27436 32376 27488 32385
rect 28172 32419 28224 32428
rect 28172 32385 28181 32419
rect 28181 32385 28215 32419
rect 28215 32385 28224 32419
rect 28172 32376 28224 32385
rect 29552 32376 29604 32428
rect 18604 32172 18656 32224
rect 19432 32172 19484 32224
rect 20168 32172 20220 32224
rect 21916 32172 21968 32224
rect 24400 32172 24452 32224
rect 25320 32215 25372 32224
rect 25320 32181 25329 32215
rect 25329 32181 25363 32215
rect 25363 32181 25372 32215
rect 28448 32240 28500 32292
rect 30380 32419 30432 32428
rect 30380 32385 30389 32419
rect 30389 32385 30423 32419
rect 30423 32385 30432 32419
rect 31300 32419 31352 32428
rect 30380 32376 30432 32385
rect 31300 32385 31309 32419
rect 31309 32385 31343 32419
rect 31343 32385 31352 32419
rect 31300 32376 31352 32385
rect 31484 32419 31536 32428
rect 31484 32385 31493 32419
rect 31493 32385 31527 32419
rect 31527 32385 31536 32419
rect 31484 32376 31536 32385
rect 32496 32512 32548 32564
rect 33784 32555 33836 32564
rect 32220 32376 32272 32428
rect 32312 32419 32364 32428
rect 32312 32385 32321 32419
rect 32321 32385 32355 32419
rect 32355 32385 32364 32419
rect 32312 32376 32364 32385
rect 30564 32308 30616 32360
rect 30932 32308 30984 32360
rect 26976 32215 27028 32224
rect 25320 32172 25372 32181
rect 26976 32181 26985 32215
rect 26985 32181 27019 32215
rect 27019 32181 27028 32215
rect 26976 32172 27028 32181
rect 28908 32172 28960 32224
rect 31024 32240 31076 32292
rect 30196 32172 30248 32224
rect 31116 32215 31168 32224
rect 31116 32181 31125 32215
rect 31125 32181 31159 32215
rect 31159 32181 31168 32215
rect 31116 32172 31168 32181
rect 31576 32351 31628 32360
rect 31576 32317 31585 32351
rect 31585 32317 31619 32351
rect 31619 32317 31628 32351
rect 31576 32308 31628 32317
rect 31760 32308 31812 32360
rect 32680 32444 32732 32496
rect 33784 32521 33793 32555
rect 33793 32521 33827 32555
rect 33827 32521 33836 32555
rect 33784 32512 33836 32521
rect 33508 32444 33560 32496
rect 33876 32444 33928 32496
rect 31484 32240 31536 32292
rect 34704 32240 34756 32292
rect 31760 32172 31812 32224
rect 33324 32215 33376 32224
rect 33324 32181 33333 32215
rect 33333 32181 33367 32215
rect 33367 32181 33376 32215
rect 33324 32172 33376 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 15292 32011 15344 32020
rect 15292 31977 15301 32011
rect 15301 31977 15335 32011
rect 15335 31977 15344 32011
rect 15292 31968 15344 31977
rect 16304 32011 16356 32020
rect 16304 31977 16313 32011
rect 16313 31977 16347 32011
rect 16347 31977 16356 32011
rect 16304 31968 16356 31977
rect 17316 31968 17368 32020
rect 20352 31968 20404 32020
rect 23204 32011 23256 32020
rect 23204 31977 23213 32011
rect 23213 31977 23247 32011
rect 23247 31977 23256 32011
rect 23204 31968 23256 31977
rect 25320 31968 25372 32020
rect 25688 31968 25740 32020
rect 26516 31968 26568 32020
rect 26976 31968 27028 32020
rect 32956 31968 33008 32020
rect 33508 32011 33560 32020
rect 33508 31977 33517 32011
rect 33517 31977 33551 32011
rect 33551 31977 33560 32011
rect 33508 31968 33560 31977
rect 15660 31832 15712 31884
rect 18788 31900 18840 31952
rect 21088 31900 21140 31952
rect 16212 31832 16264 31884
rect 18604 31832 18656 31884
rect 25044 31900 25096 31952
rect 22284 31875 22336 31884
rect 22284 31841 22293 31875
rect 22293 31841 22327 31875
rect 22327 31841 22336 31875
rect 22284 31832 22336 31841
rect 24584 31832 24636 31884
rect 27528 31832 27580 31884
rect 15476 31807 15528 31816
rect 15476 31773 15485 31807
rect 15485 31773 15519 31807
rect 15519 31773 15528 31807
rect 15476 31764 15528 31773
rect 16764 31807 16816 31816
rect 16028 31696 16080 31748
rect 15936 31628 15988 31680
rect 16764 31773 16773 31807
rect 16773 31773 16807 31807
rect 16807 31773 16816 31807
rect 16764 31764 16816 31773
rect 16856 31807 16908 31816
rect 16856 31773 16865 31807
rect 16865 31773 16899 31807
rect 16899 31773 16908 31807
rect 19432 31807 19484 31816
rect 16856 31764 16908 31773
rect 17040 31696 17092 31748
rect 19432 31773 19441 31807
rect 19441 31773 19475 31807
rect 19475 31773 19484 31807
rect 19432 31764 19484 31773
rect 21088 31807 21140 31816
rect 20168 31696 20220 31748
rect 21088 31773 21097 31807
rect 21097 31773 21131 31807
rect 21131 31773 21140 31807
rect 21088 31764 21140 31773
rect 21916 31807 21968 31816
rect 21916 31773 21925 31807
rect 21925 31773 21959 31807
rect 21959 31773 21968 31807
rect 21916 31764 21968 31773
rect 26148 31807 26200 31816
rect 26148 31773 26157 31807
rect 26157 31773 26191 31807
rect 26191 31773 26200 31807
rect 26148 31764 26200 31773
rect 23756 31739 23808 31748
rect 23756 31705 23765 31739
rect 23765 31705 23799 31739
rect 23799 31705 23808 31739
rect 23756 31696 23808 31705
rect 24400 31696 24452 31748
rect 25964 31696 26016 31748
rect 28172 31764 28224 31816
rect 28448 31807 28500 31816
rect 28448 31773 28457 31807
rect 28457 31773 28491 31807
rect 28491 31773 28500 31807
rect 28448 31764 28500 31773
rect 29092 31900 29144 31952
rect 29552 31875 29604 31884
rect 29552 31841 29561 31875
rect 29561 31841 29595 31875
rect 29595 31841 29604 31875
rect 29552 31832 29604 31841
rect 30564 31832 30616 31884
rect 18052 31628 18104 31680
rect 18236 31628 18288 31680
rect 19432 31628 19484 31680
rect 20720 31628 20772 31680
rect 21824 31628 21876 31680
rect 21916 31628 21968 31680
rect 23388 31628 23440 31680
rect 23480 31628 23532 31680
rect 23848 31628 23900 31680
rect 25688 31628 25740 31680
rect 28540 31696 28592 31748
rect 30196 31764 30248 31816
rect 31576 31900 31628 31952
rect 32588 31900 32640 31952
rect 35624 31968 35676 32020
rect 30932 31832 30984 31884
rect 31392 31807 31444 31816
rect 31392 31773 31401 31807
rect 31401 31773 31435 31807
rect 31435 31773 31444 31807
rect 31392 31764 31444 31773
rect 32220 31807 32272 31816
rect 31484 31696 31536 31748
rect 32220 31773 32229 31807
rect 32229 31773 32263 31807
rect 32263 31773 32272 31807
rect 32220 31764 32272 31773
rect 32312 31807 32364 31816
rect 32312 31773 32321 31807
rect 32321 31773 32355 31807
rect 32355 31773 32364 31807
rect 33048 31832 33100 31884
rect 33232 31832 33284 31884
rect 34152 31900 34204 31952
rect 34704 31900 34756 31952
rect 36084 31900 36136 31952
rect 35532 31832 35584 31884
rect 32312 31764 32364 31773
rect 32588 31807 32640 31816
rect 32588 31773 32597 31807
rect 32597 31773 32631 31807
rect 32631 31773 32640 31807
rect 32588 31764 32640 31773
rect 32956 31764 33008 31816
rect 33416 31764 33468 31816
rect 31852 31696 31904 31748
rect 34152 31807 34204 31816
rect 34152 31773 34161 31807
rect 34161 31773 34195 31807
rect 34195 31773 34204 31807
rect 34152 31764 34204 31773
rect 34704 31807 34756 31816
rect 34704 31773 34713 31807
rect 34713 31773 34747 31807
rect 34747 31773 34756 31807
rect 34704 31764 34756 31773
rect 34060 31696 34112 31748
rect 28724 31628 28776 31680
rect 31576 31628 31628 31680
rect 32036 31671 32088 31680
rect 32036 31637 32045 31671
rect 32045 31637 32079 31671
rect 32079 31637 32088 31671
rect 32036 31628 32088 31637
rect 34520 31628 34572 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 15476 31424 15528 31476
rect 16028 31424 16080 31476
rect 16856 31467 16908 31476
rect 16856 31433 16865 31467
rect 16865 31433 16899 31467
rect 16899 31433 16908 31467
rect 16856 31424 16908 31433
rect 18328 31467 18380 31476
rect 18328 31433 18337 31467
rect 18337 31433 18371 31467
rect 18371 31433 18380 31467
rect 18328 31424 18380 31433
rect 18788 31467 18840 31476
rect 18788 31433 18797 31467
rect 18797 31433 18831 31467
rect 18831 31433 18840 31467
rect 18788 31424 18840 31433
rect 19248 31424 19300 31476
rect 19340 31424 19392 31476
rect 15292 31331 15344 31340
rect 15292 31297 15301 31331
rect 15301 31297 15335 31331
rect 15335 31297 15344 31331
rect 15292 31288 15344 31297
rect 16028 31288 16080 31340
rect 16856 31288 16908 31340
rect 17040 31331 17092 31340
rect 17040 31297 17049 31331
rect 17049 31297 17083 31331
rect 17083 31297 17092 31331
rect 17040 31288 17092 31297
rect 15844 31220 15896 31272
rect 17868 31288 17920 31340
rect 19432 31356 19484 31408
rect 20260 31424 20312 31476
rect 24584 31467 24636 31476
rect 24584 31433 24593 31467
rect 24593 31433 24627 31467
rect 24627 31433 24636 31467
rect 24584 31424 24636 31433
rect 26792 31424 26844 31476
rect 18512 31288 18564 31340
rect 18972 31331 19024 31340
rect 18972 31297 18981 31331
rect 18981 31297 19015 31331
rect 19015 31297 19024 31331
rect 18972 31288 19024 31297
rect 17960 31220 18012 31272
rect 15200 31152 15252 31204
rect 18052 31152 18104 31204
rect 19156 31288 19208 31340
rect 20076 31331 20128 31340
rect 20076 31297 20085 31331
rect 20085 31297 20119 31331
rect 20119 31297 20128 31331
rect 20076 31288 20128 31297
rect 21180 31331 21232 31340
rect 20168 31263 20220 31272
rect 20168 31229 20177 31263
rect 20177 31229 20211 31263
rect 20211 31229 20220 31263
rect 20168 31220 20220 31229
rect 20260 31152 20312 31204
rect 20720 31152 20772 31204
rect 21180 31297 21189 31331
rect 21189 31297 21223 31331
rect 21223 31297 21232 31331
rect 21180 31288 21232 31297
rect 21824 31288 21876 31340
rect 23112 31288 23164 31340
rect 24676 31356 24728 31408
rect 26056 31356 26108 31408
rect 24032 31331 24084 31340
rect 24032 31297 24041 31331
rect 24041 31297 24075 31331
rect 24075 31297 24084 31331
rect 24032 31288 24084 31297
rect 21088 31220 21140 31272
rect 22008 31263 22060 31272
rect 22008 31229 22017 31263
rect 22017 31229 22051 31263
rect 22051 31229 22060 31263
rect 22008 31220 22060 31229
rect 21456 31152 21508 31204
rect 21916 31152 21968 31204
rect 22744 31220 22796 31272
rect 24952 31288 25004 31340
rect 25780 31288 25832 31340
rect 26424 31288 26476 31340
rect 26792 31288 26844 31340
rect 27528 31424 27580 31476
rect 30564 31424 30616 31476
rect 33140 31467 33192 31476
rect 27252 31399 27304 31408
rect 27252 31365 27261 31399
rect 27261 31365 27295 31399
rect 27295 31365 27304 31399
rect 27252 31356 27304 31365
rect 30472 31356 30524 31408
rect 26332 31152 26384 31204
rect 26608 31152 26660 31204
rect 28540 31288 28592 31340
rect 29092 31331 29144 31340
rect 15292 31084 15344 31136
rect 16948 31084 17000 31136
rect 18144 31127 18196 31136
rect 18144 31093 18153 31127
rect 18153 31093 18187 31127
rect 18187 31093 18196 31127
rect 18144 31084 18196 31093
rect 19984 31084 20036 31136
rect 23204 31084 23256 31136
rect 23940 31127 23992 31136
rect 23940 31093 23949 31127
rect 23949 31093 23983 31127
rect 23983 31093 23992 31127
rect 23940 31084 23992 31093
rect 27252 31084 27304 31136
rect 28080 31127 28132 31136
rect 28080 31093 28089 31127
rect 28089 31093 28123 31127
rect 28123 31093 28132 31127
rect 28080 31084 28132 31093
rect 28264 31152 28316 31204
rect 29092 31297 29101 31331
rect 29101 31297 29135 31331
rect 29135 31297 29144 31331
rect 29092 31288 29144 31297
rect 29828 31288 29880 31340
rect 30932 31331 30984 31340
rect 29552 31220 29604 31272
rect 30472 31220 30524 31272
rect 29828 31152 29880 31204
rect 30932 31297 30941 31331
rect 30941 31297 30975 31331
rect 30975 31297 30984 31331
rect 30932 31288 30984 31297
rect 33140 31433 33149 31467
rect 33149 31433 33183 31467
rect 33183 31433 33192 31467
rect 33140 31424 33192 31433
rect 31300 31356 31352 31408
rect 31852 31288 31904 31340
rect 32128 31288 32180 31340
rect 34520 31331 34572 31340
rect 30104 31127 30156 31136
rect 30104 31093 30113 31127
rect 30113 31093 30147 31127
rect 30147 31093 30156 31127
rect 30104 31084 30156 31093
rect 30472 31084 30524 31136
rect 32036 31220 32088 31272
rect 32588 31220 32640 31272
rect 32864 31220 32916 31272
rect 34520 31297 34529 31331
rect 34529 31297 34563 31331
rect 34563 31297 34572 31331
rect 34520 31288 34572 31297
rect 35532 31331 35584 31340
rect 35532 31297 35541 31331
rect 35541 31297 35575 31331
rect 35575 31297 35584 31331
rect 35532 31288 35584 31297
rect 34612 31263 34664 31272
rect 34612 31229 34621 31263
rect 34621 31229 34655 31263
rect 34655 31229 34664 31263
rect 34612 31220 34664 31229
rect 31208 31152 31260 31204
rect 35992 31152 36044 31204
rect 31484 31084 31536 31136
rect 31668 31084 31720 31136
rect 32680 31084 32732 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 15200 30923 15252 30932
rect 15200 30889 15209 30923
rect 15209 30889 15243 30923
rect 15243 30889 15252 30923
rect 15200 30880 15252 30889
rect 16764 30880 16816 30932
rect 16028 30744 16080 30796
rect 15660 30719 15712 30728
rect 15660 30685 15669 30719
rect 15669 30685 15703 30719
rect 15703 30685 15712 30719
rect 15660 30676 15712 30685
rect 15936 30676 15988 30728
rect 16580 30719 16632 30728
rect 16580 30685 16589 30719
rect 16589 30685 16623 30719
rect 16623 30685 16632 30719
rect 16580 30676 16632 30685
rect 15844 30540 15896 30592
rect 16764 30651 16816 30660
rect 16764 30617 16773 30651
rect 16773 30617 16807 30651
rect 16807 30617 16816 30651
rect 17592 30676 17644 30728
rect 18236 30880 18288 30932
rect 20076 30880 20128 30932
rect 21088 30880 21140 30932
rect 23112 30880 23164 30932
rect 29736 30923 29788 30932
rect 17960 30812 18012 30864
rect 18144 30855 18196 30864
rect 18144 30821 18153 30855
rect 18153 30821 18187 30855
rect 18187 30821 18196 30855
rect 18144 30812 18196 30821
rect 23020 30812 23072 30864
rect 23480 30855 23532 30864
rect 23480 30821 23489 30855
rect 23489 30821 23523 30855
rect 23523 30821 23532 30855
rect 23480 30812 23532 30821
rect 24952 30812 25004 30864
rect 23204 30787 23256 30796
rect 16764 30608 16816 30617
rect 17040 30540 17092 30592
rect 17776 30540 17828 30592
rect 18052 30676 18104 30728
rect 18328 30676 18380 30728
rect 19524 30676 19576 30728
rect 19340 30608 19392 30660
rect 21456 30719 21508 30728
rect 21456 30685 21465 30719
rect 21465 30685 21499 30719
rect 21499 30685 21508 30719
rect 21456 30676 21508 30685
rect 23204 30753 23213 30787
rect 23213 30753 23247 30787
rect 23247 30753 23256 30787
rect 23204 30744 23256 30753
rect 22192 30719 22244 30728
rect 21272 30608 21324 30660
rect 22192 30685 22201 30719
rect 22201 30685 22235 30719
rect 22235 30685 22244 30719
rect 22192 30676 22244 30685
rect 22376 30719 22428 30728
rect 22376 30685 22385 30719
rect 22385 30685 22419 30719
rect 22419 30685 22428 30719
rect 22376 30676 22428 30685
rect 23940 30676 23992 30728
rect 26700 30744 26752 30796
rect 26240 30719 26292 30728
rect 26240 30685 26249 30719
rect 26249 30685 26283 30719
rect 26283 30685 26292 30719
rect 26240 30676 26292 30685
rect 28908 30812 28960 30864
rect 28080 30744 28132 30796
rect 28356 30744 28408 30796
rect 29736 30889 29745 30923
rect 29745 30889 29779 30923
rect 29779 30889 29788 30923
rect 29736 30880 29788 30889
rect 30380 30880 30432 30932
rect 31024 30880 31076 30932
rect 31484 30923 31536 30932
rect 31484 30889 31493 30923
rect 31493 30889 31527 30923
rect 31527 30889 31536 30923
rect 31484 30880 31536 30889
rect 31576 30923 31628 30932
rect 31576 30889 31585 30923
rect 31585 30889 31619 30923
rect 31619 30889 31628 30923
rect 31576 30880 31628 30889
rect 32680 30923 32732 30932
rect 30104 30812 30156 30864
rect 31852 30812 31904 30864
rect 32680 30889 32689 30923
rect 32689 30889 32723 30923
rect 32723 30889 32732 30923
rect 32680 30880 32732 30889
rect 33968 30880 34020 30932
rect 31576 30744 31628 30796
rect 33324 30812 33376 30864
rect 35992 30787 36044 30796
rect 22836 30608 22888 30660
rect 25228 30608 25280 30660
rect 26332 30608 26384 30660
rect 27252 30719 27304 30728
rect 27252 30685 27261 30719
rect 27261 30685 27295 30719
rect 27295 30685 27304 30719
rect 27252 30676 27304 30685
rect 28540 30676 28592 30728
rect 29000 30676 29052 30728
rect 31116 30676 31168 30728
rect 30932 30608 30984 30660
rect 31392 30608 31444 30660
rect 18052 30540 18104 30592
rect 18604 30540 18656 30592
rect 21640 30583 21692 30592
rect 21640 30549 21649 30583
rect 21649 30549 21683 30583
rect 21683 30549 21692 30583
rect 21640 30540 21692 30549
rect 21732 30540 21784 30592
rect 25412 30583 25464 30592
rect 25412 30549 25421 30583
rect 25421 30549 25455 30583
rect 25455 30549 25464 30583
rect 25412 30540 25464 30549
rect 26148 30583 26200 30592
rect 26148 30549 26157 30583
rect 26157 30549 26191 30583
rect 26191 30549 26200 30583
rect 26148 30540 26200 30549
rect 27344 30540 27396 30592
rect 28816 30540 28868 30592
rect 29460 30540 29512 30592
rect 30288 30540 30340 30592
rect 35992 30753 36001 30787
rect 36001 30753 36035 30787
rect 36035 30753 36044 30787
rect 35992 30744 36044 30753
rect 32588 30676 32640 30728
rect 33600 30719 33652 30728
rect 32128 30540 32180 30592
rect 32772 30608 32824 30660
rect 33600 30685 33609 30719
rect 33609 30685 33643 30719
rect 33643 30685 33652 30719
rect 33600 30676 33652 30685
rect 35072 30719 35124 30728
rect 35072 30685 35081 30719
rect 35081 30685 35115 30719
rect 35115 30685 35124 30719
rect 35072 30676 35124 30685
rect 35624 30676 35676 30728
rect 35900 30719 35952 30728
rect 35900 30685 35909 30719
rect 35909 30685 35943 30719
rect 35943 30685 35952 30719
rect 35900 30676 35952 30685
rect 34060 30608 34112 30660
rect 36176 30540 36228 30592
rect 37188 30540 37240 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 15660 30268 15712 30320
rect 15936 30336 15988 30388
rect 17868 30336 17920 30388
rect 18328 30336 18380 30388
rect 18512 30379 18564 30388
rect 18512 30345 18521 30379
rect 18521 30345 18555 30379
rect 18555 30345 18564 30379
rect 18512 30336 18564 30345
rect 21456 30336 21508 30388
rect 22100 30336 22152 30388
rect 22744 30336 22796 30388
rect 23204 30336 23256 30388
rect 23848 30336 23900 30388
rect 26240 30336 26292 30388
rect 28540 30336 28592 30388
rect 30380 30336 30432 30388
rect 31300 30336 31352 30388
rect 35072 30336 35124 30388
rect 20812 30311 20864 30320
rect 20812 30277 20821 30311
rect 20821 30277 20855 30311
rect 20855 30277 20864 30311
rect 20812 30268 20864 30277
rect 21640 30268 21692 30320
rect 24124 30268 24176 30320
rect 15844 30243 15896 30252
rect 15844 30209 15853 30243
rect 15853 30209 15887 30243
rect 15887 30209 15896 30243
rect 15844 30200 15896 30209
rect 16580 30200 16632 30252
rect 17040 30243 17092 30252
rect 17040 30209 17049 30243
rect 17049 30209 17083 30243
rect 17083 30209 17092 30243
rect 17040 30200 17092 30209
rect 16764 30132 16816 30184
rect 17592 30200 17644 30252
rect 19248 30243 19300 30252
rect 19248 30209 19257 30243
rect 19257 30209 19291 30243
rect 19291 30209 19300 30243
rect 19248 30200 19300 30209
rect 19432 30243 19484 30252
rect 19432 30209 19441 30243
rect 19441 30209 19475 30243
rect 19475 30209 19484 30243
rect 19432 30200 19484 30209
rect 17776 30175 17828 30184
rect 17776 30141 17785 30175
rect 17785 30141 17819 30175
rect 17819 30141 17828 30175
rect 17776 30132 17828 30141
rect 19156 30175 19208 30184
rect 19156 30141 19165 30175
rect 19165 30141 19199 30175
rect 19199 30141 19208 30175
rect 19156 30132 19208 30141
rect 20352 30200 20404 30252
rect 21364 30200 21416 30252
rect 21824 30243 21876 30252
rect 21824 30209 21833 30243
rect 21833 30209 21867 30243
rect 21867 30209 21876 30243
rect 21824 30200 21876 30209
rect 22008 30243 22060 30252
rect 22008 30209 22017 30243
rect 22017 30209 22051 30243
rect 22051 30209 22060 30243
rect 22008 30200 22060 30209
rect 22744 30200 22796 30252
rect 24584 30200 24636 30252
rect 25228 30243 25280 30252
rect 25228 30209 25237 30243
rect 25237 30209 25271 30243
rect 25271 30209 25280 30243
rect 25228 30200 25280 30209
rect 25320 30200 25372 30252
rect 26148 30200 26200 30252
rect 26516 30200 26568 30252
rect 28080 30268 28132 30320
rect 29092 30268 29144 30320
rect 20260 30175 20312 30184
rect 20260 30141 20269 30175
rect 20269 30141 20303 30175
rect 20303 30141 20312 30175
rect 20260 30132 20312 30141
rect 23112 30132 23164 30184
rect 25044 30132 25096 30184
rect 16948 30064 17000 30116
rect 22468 30064 22520 30116
rect 23572 30064 23624 30116
rect 24124 30064 24176 30116
rect 24768 30064 24820 30116
rect 24952 30064 25004 30116
rect 27528 30132 27580 30184
rect 27620 30209 27629 30218
rect 27629 30209 27663 30218
rect 27663 30209 27672 30218
rect 27620 30166 27672 30209
rect 27804 30243 27856 30252
rect 27804 30209 27813 30243
rect 27813 30209 27847 30243
rect 27847 30209 27856 30243
rect 27804 30200 27856 30209
rect 28448 30200 28500 30252
rect 29736 30200 29788 30252
rect 28172 30132 28224 30184
rect 28264 30132 28316 30184
rect 31944 30200 31996 30252
rect 32220 30268 32272 30320
rect 32956 30268 33008 30320
rect 35624 30268 35676 30320
rect 29920 30132 29972 30184
rect 30288 30175 30340 30184
rect 30288 30141 30297 30175
rect 30297 30141 30331 30175
rect 30331 30141 30340 30175
rect 30288 30132 30340 30141
rect 30472 30132 30524 30184
rect 32496 30200 32548 30252
rect 33048 30243 33100 30252
rect 33048 30209 33057 30243
rect 33057 30209 33091 30243
rect 33091 30209 33100 30243
rect 33048 30200 33100 30209
rect 34152 30243 34204 30252
rect 34152 30209 34161 30243
rect 34161 30209 34195 30243
rect 34195 30209 34204 30243
rect 34152 30200 34204 30209
rect 36268 30243 36320 30252
rect 36268 30209 36277 30243
rect 36277 30209 36311 30243
rect 36311 30209 36320 30243
rect 36268 30200 36320 30209
rect 37924 30200 37976 30252
rect 36176 30175 36228 30184
rect 36176 30141 36185 30175
rect 36185 30141 36219 30175
rect 36219 30141 36228 30175
rect 36176 30132 36228 30141
rect 37372 30175 37424 30184
rect 37372 30141 37381 30175
rect 37381 30141 37415 30175
rect 37415 30141 37424 30175
rect 37372 30132 37424 30141
rect 16580 29996 16632 30048
rect 17776 29996 17828 30048
rect 22652 29996 22704 30048
rect 22836 30039 22888 30048
rect 22836 30005 22845 30039
rect 22845 30005 22879 30039
rect 22879 30005 22888 30039
rect 22836 29996 22888 30005
rect 22928 29996 22980 30048
rect 28080 29996 28132 30048
rect 28632 29996 28684 30048
rect 30932 29996 30984 30048
rect 32312 29996 32364 30048
rect 33968 29996 34020 30048
rect 34796 30064 34848 30116
rect 37832 30107 37884 30116
rect 37832 30073 37841 30107
rect 37841 30073 37875 30107
rect 37875 30073 37884 30107
rect 37832 30064 37884 30073
rect 35900 29996 35952 30048
rect 36544 30039 36596 30048
rect 36544 30005 36553 30039
rect 36553 30005 36587 30039
rect 36587 30005 36596 30039
rect 36544 29996 36596 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 17040 29792 17092 29844
rect 18052 29835 18104 29844
rect 18052 29801 18061 29835
rect 18061 29801 18095 29835
rect 18095 29801 18104 29835
rect 18052 29792 18104 29801
rect 19340 29792 19392 29844
rect 20076 29792 20128 29844
rect 21272 29835 21324 29844
rect 21272 29801 21281 29835
rect 21281 29801 21315 29835
rect 21315 29801 21324 29835
rect 21272 29792 21324 29801
rect 22836 29792 22888 29844
rect 23020 29792 23072 29844
rect 22468 29724 22520 29776
rect 25228 29792 25280 29844
rect 16028 29656 16080 29708
rect 17408 29656 17460 29708
rect 16580 29588 16632 29640
rect 17960 29631 18012 29640
rect 17960 29597 17969 29631
rect 17969 29597 18003 29631
rect 18003 29597 18012 29631
rect 17960 29588 18012 29597
rect 18236 29588 18288 29640
rect 21088 29631 21140 29640
rect 15476 29520 15528 29572
rect 15844 29520 15896 29572
rect 16120 29520 16172 29572
rect 20260 29520 20312 29572
rect 21088 29597 21097 29631
rect 21097 29597 21131 29631
rect 21131 29597 21140 29631
rect 21088 29588 21140 29597
rect 22744 29588 22796 29640
rect 23388 29631 23440 29640
rect 23388 29597 23397 29631
rect 23397 29597 23431 29631
rect 23431 29597 23440 29631
rect 23388 29588 23440 29597
rect 24216 29656 24268 29708
rect 22100 29520 22152 29572
rect 19984 29495 20036 29504
rect 19984 29461 20009 29495
rect 20009 29461 20036 29495
rect 20168 29495 20220 29504
rect 19984 29452 20036 29461
rect 20168 29461 20177 29495
rect 20177 29461 20211 29495
rect 20211 29461 20220 29495
rect 20168 29452 20220 29461
rect 22468 29452 22520 29504
rect 24124 29520 24176 29572
rect 25044 29724 25096 29776
rect 25688 29767 25740 29776
rect 24676 29699 24728 29708
rect 24676 29665 24685 29699
rect 24685 29665 24719 29699
rect 24719 29665 24728 29699
rect 24676 29656 24728 29665
rect 24768 29588 24820 29640
rect 25228 29656 25280 29708
rect 25412 29699 25464 29708
rect 25412 29665 25421 29699
rect 25421 29665 25455 29699
rect 25455 29665 25464 29699
rect 25412 29656 25464 29665
rect 25688 29733 25697 29767
rect 25697 29733 25731 29767
rect 25731 29733 25740 29767
rect 25688 29724 25740 29733
rect 29000 29792 29052 29844
rect 29368 29792 29420 29844
rect 34704 29792 34756 29844
rect 37372 29792 37424 29844
rect 25320 29631 25372 29640
rect 25320 29597 25329 29631
rect 25329 29597 25363 29631
rect 25363 29597 25372 29631
rect 25320 29588 25372 29597
rect 28908 29656 28960 29708
rect 29092 29656 29144 29708
rect 33600 29724 33652 29776
rect 34152 29724 34204 29776
rect 30656 29656 30708 29708
rect 31852 29699 31904 29708
rect 28080 29588 28132 29640
rect 26148 29563 26200 29572
rect 26148 29529 26157 29563
rect 26157 29529 26191 29563
rect 26191 29529 26200 29563
rect 26148 29520 26200 29529
rect 29184 29520 29236 29572
rect 30012 29563 30064 29572
rect 30012 29529 30021 29563
rect 30021 29529 30055 29563
rect 30055 29529 30064 29563
rect 30012 29520 30064 29529
rect 31208 29588 31260 29640
rect 31852 29665 31861 29699
rect 31861 29665 31895 29699
rect 31895 29665 31904 29699
rect 31852 29656 31904 29665
rect 32220 29656 32272 29708
rect 32864 29656 32916 29708
rect 33232 29699 33284 29708
rect 33232 29665 33241 29699
rect 33241 29665 33275 29699
rect 33275 29665 33284 29699
rect 33232 29656 33284 29665
rect 36268 29724 36320 29776
rect 32496 29588 32548 29640
rect 34796 29656 34848 29708
rect 33968 29588 34020 29640
rect 34520 29588 34572 29640
rect 34704 29631 34756 29640
rect 34704 29597 34713 29631
rect 34713 29597 34747 29631
rect 34747 29597 34756 29631
rect 34704 29588 34756 29597
rect 34980 29588 35032 29640
rect 23480 29452 23532 29504
rect 23756 29452 23808 29504
rect 24032 29452 24084 29504
rect 24584 29452 24636 29504
rect 27252 29452 27304 29504
rect 28172 29452 28224 29504
rect 29276 29452 29328 29504
rect 29920 29452 29972 29504
rect 30104 29452 30156 29504
rect 33784 29520 33836 29572
rect 35624 29588 35676 29640
rect 36176 29588 36228 29640
rect 36268 29563 36320 29572
rect 36268 29529 36277 29563
rect 36277 29529 36311 29563
rect 36311 29529 36320 29563
rect 36268 29520 36320 29529
rect 32220 29452 32272 29504
rect 32956 29452 33008 29504
rect 34888 29452 34940 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 17408 29291 17460 29300
rect 17408 29257 17417 29291
rect 17417 29257 17451 29291
rect 17451 29257 17460 29291
rect 17408 29248 17460 29257
rect 17776 29291 17828 29300
rect 17776 29257 17785 29291
rect 17785 29257 17819 29291
rect 17819 29257 17828 29291
rect 17776 29248 17828 29257
rect 15844 29180 15896 29232
rect 16948 29223 17000 29232
rect 16948 29189 16957 29223
rect 16957 29189 16991 29223
rect 16991 29189 17000 29223
rect 16948 29180 17000 29189
rect 16120 29155 16172 29164
rect 16120 29121 16129 29155
rect 16129 29121 16163 29155
rect 16163 29121 16172 29155
rect 16120 29112 16172 29121
rect 17592 29155 17644 29164
rect 17592 29121 17601 29155
rect 17601 29121 17635 29155
rect 17635 29121 17644 29155
rect 17592 29112 17644 29121
rect 17868 29155 17920 29164
rect 17868 29121 17877 29155
rect 17877 29121 17911 29155
rect 17911 29121 17920 29155
rect 17868 29112 17920 29121
rect 19984 29180 20036 29232
rect 22192 29248 22244 29300
rect 21088 29180 21140 29232
rect 18512 29155 18564 29164
rect 18236 29044 18288 29096
rect 18512 29121 18521 29155
rect 18521 29121 18555 29155
rect 18555 29121 18564 29155
rect 18512 29112 18564 29121
rect 19708 29155 19760 29164
rect 18604 29044 18656 29096
rect 19708 29121 19717 29155
rect 19717 29121 19751 29155
rect 19751 29121 19760 29155
rect 19708 29112 19760 29121
rect 20076 29112 20128 29164
rect 20260 29155 20312 29164
rect 20260 29121 20269 29155
rect 20269 29121 20303 29155
rect 20303 29121 20312 29155
rect 20260 29112 20312 29121
rect 20352 29112 20404 29164
rect 20904 29112 20956 29164
rect 21916 29112 21968 29164
rect 23020 29112 23072 29164
rect 23848 29155 23900 29164
rect 23848 29121 23857 29155
rect 23857 29121 23891 29155
rect 23891 29121 23900 29155
rect 23848 29112 23900 29121
rect 24768 29248 24820 29300
rect 24109 29155 24161 29164
rect 24109 29121 24126 29155
rect 24126 29121 24161 29155
rect 24109 29112 24161 29121
rect 24216 29155 24268 29164
rect 26148 29248 26200 29300
rect 27620 29248 27672 29300
rect 28080 29291 28132 29300
rect 28080 29257 28089 29291
rect 28089 29257 28123 29291
rect 28123 29257 28132 29291
rect 28080 29248 28132 29257
rect 28724 29291 28776 29300
rect 25228 29180 25280 29232
rect 24216 29121 24235 29155
rect 24235 29121 24268 29155
rect 24216 29112 24268 29121
rect 21732 29044 21784 29096
rect 25044 29155 25096 29164
rect 25044 29121 25053 29155
rect 25053 29121 25087 29155
rect 25087 29121 25096 29155
rect 25044 29112 25096 29121
rect 20720 28976 20772 29028
rect 24584 29044 24636 29096
rect 24400 28976 24452 29028
rect 26516 29112 26568 29164
rect 27160 29180 27212 29232
rect 28724 29257 28749 29291
rect 28749 29257 28776 29291
rect 28724 29248 28776 29257
rect 28540 29223 28592 29232
rect 28540 29189 28549 29223
rect 28549 29189 28583 29223
rect 28583 29189 28592 29223
rect 30012 29248 30064 29300
rect 31944 29248 31996 29300
rect 32312 29291 32364 29300
rect 32312 29257 32337 29291
rect 32337 29257 32364 29291
rect 32312 29248 32364 29257
rect 28540 29180 28592 29189
rect 28908 29180 28960 29232
rect 29092 29180 29144 29232
rect 26608 29044 26660 29096
rect 29276 29112 29328 29164
rect 29460 29155 29512 29164
rect 29460 29121 29469 29155
rect 29469 29121 29503 29155
rect 29503 29121 29512 29155
rect 29460 29112 29512 29121
rect 27252 29044 27304 29096
rect 27712 28976 27764 29028
rect 29368 29044 29420 29096
rect 32036 29180 32088 29232
rect 32680 29248 32732 29300
rect 33048 29248 33100 29300
rect 33232 29291 33284 29300
rect 33232 29257 33241 29291
rect 33241 29257 33275 29291
rect 33275 29257 33284 29291
rect 33232 29248 33284 29257
rect 34336 29248 34388 29300
rect 34980 29248 35032 29300
rect 37924 29291 37976 29300
rect 37924 29257 37933 29291
rect 37933 29257 37967 29291
rect 37967 29257 37976 29291
rect 37924 29248 37976 29257
rect 34796 29180 34848 29232
rect 36544 29180 36596 29232
rect 29644 29044 29696 29096
rect 30380 29112 30432 29164
rect 30656 29155 30708 29164
rect 30656 29121 30665 29155
rect 30665 29121 30699 29155
rect 30699 29121 30708 29155
rect 30656 29112 30708 29121
rect 31208 29155 31260 29164
rect 31208 29121 31217 29155
rect 31217 29121 31251 29155
rect 31251 29121 31260 29155
rect 31208 29112 31260 29121
rect 32956 29155 33008 29164
rect 32956 29121 32965 29155
rect 32965 29121 32999 29155
rect 32999 29121 33008 29155
rect 32956 29112 33008 29121
rect 33876 29155 33928 29164
rect 33876 29121 33885 29155
rect 33885 29121 33919 29155
rect 33919 29121 33928 29155
rect 33876 29112 33928 29121
rect 34704 29155 34756 29164
rect 34704 29121 34713 29155
rect 34713 29121 34747 29155
rect 34747 29121 34756 29155
rect 34704 29112 34756 29121
rect 34888 29112 34940 29164
rect 30104 29044 30156 29096
rect 33232 29087 33284 29096
rect 33232 29053 33241 29087
rect 33241 29053 33275 29087
rect 33275 29053 33284 29087
rect 33232 29044 33284 29053
rect 33968 29087 34020 29096
rect 33968 29053 33977 29087
rect 33977 29053 34011 29087
rect 34011 29053 34020 29087
rect 33968 29044 34020 29053
rect 34520 29044 34572 29096
rect 28448 28976 28500 29028
rect 30564 29019 30616 29028
rect 18420 28951 18472 28960
rect 18420 28917 18429 28951
rect 18429 28917 18463 28951
rect 18463 28917 18472 28951
rect 18420 28908 18472 28917
rect 19248 28908 19300 28960
rect 20260 28908 20312 28960
rect 20536 28908 20588 28960
rect 20904 28908 20956 28960
rect 24584 28908 24636 28960
rect 24952 28908 25004 28960
rect 25872 28908 25924 28960
rect 29460 28908 29512 28960
rect 29736 28908 29788 28960
rect 30104 28908 30156 28960
rect 30564 28985 30573 29019
rect 30573 28985 30607 29019
rect 30607 28985 30616 29019
rect 30564 28976 30616 28985
rect 31208 28976 31260 29028
rect 32680 28976 32732 29028
rect 34152 28976 34204 29028
rect 34612 28976 34664 29028
rect 36636 29155 36688 29164
rect 36636 29121 36645 29155
rect 36645 29121 36679 29155
rect 36679 29121 36688 29155
rect 36636 29112 36688 29121
rect 35532 29087 35584 29096
rect 35532 29053 35541 29087
rect 35541 29053 35575 29087
rect 35575 29053 35584 29087
rect 37280 29087 37332 29096
rect 35532 29044 35584 29053
rect 37280 29053 37289 29087
rect 37289 29053 37323 29087
rect 37323 29053 37332 29087
rect 37280 29044 37332 29053
rect 37464 29044 37516 29096
rect 37924 28976 37976 29028
rect 31852 28908 31904 28960
rect 33048 28951 33100 28960
rect 33048 28917 33057 28951
rect 33057 28917 33091 28951
rect 33091 28917 33100 28951
rect 33048 28908 33100 28917
rect 34428 28908 34480 28960
rect 34796 28951 34848 28960
rect 34796 28917 34805 28951
rect 34805 28917 34839 28951
rect 34839 28917 34848 28951
rect 34796 28908 34848 28917
rect 35900 28951 35952 28960
rect 35900 28917 35909 28951
rect 35909 28917 35943 28951
rect 35943 28917 35952 28951
rect 35900 28908 35952 28917
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 15476 28747 15528 28756
rect 15476 28713 15485 28747
rect 15485 28713 15519 28747
rect 15519 28713 15528 28747
rect 15476 28704 15528 28713
rect 16580 28704 16632 28756
rect 17224 28704 17276 28756
rect 19156 28704 19208 28756
rect 19892 28704 19944 28756
rect 19984 28704 20036 28756
rect 19340 28636 19392 28688
rect 16028 28500 16080 28552
rect 16948 28500 17000 28552
rect 18420 28500 18472 28552
rect 16120 28475 16172 28484
rect 16120 28441 16129 28475
rect 16129 28441 16163 28475
rect 16163 28441 16172 28475
rect 16120 28432 16172 28441
rect 18328 28475 18380 28484
rect 18328 28441 18337 28475
rect 18337 28441 18371 28475
rect 18371 28441 18380 28475
rect 18328 28432 18380 28441
rect 19800 28568 19852 28620
rect 20260 28636 20312 28688
rect 22376 28704 22428 28756
rect 23848 28747 23900 28756
rect 23848 28713 23857 28747
rect 23857 28713 23891 28747
rect 23891 28713 23900 28747
rect 23848 28704 23900 28713
rect 20444 28636 20496 28688
rect 23664 28636 23716 28688
rect 27160 28704 27212 28756
rect 27620 28704 27672 28756
rect 19432 28500 19484 28552
rect 19708 28500 19760 28552
rect 19800 28432 19852 28484
rect 20444 28500 20496 28552
rect 20628 28500 20680 28552
rect 20720 28500 20772 28552
rect 21824 28543 21876 28552
rect 21824 28509 21833 28543
rect 21833 28509 21867 28543
rect 21867 28509 21876 28543
rect 21824 28500 21876 28509
rect 22008 28543 22060 28552
rect 22008 28509 22017 28543
rect 22017 28509 22051 28543
rect 22051 28509 22060 28543
rect 22008 28500 22060 28509
rect 22652 28500 22704 28552
rect 27528 28636 27580 28688
rect 27804 28568 27856 28620
rect 30380 28704 30432 28756
rect 31024 28704 31076 28756
rect 33784 28704 33836 28756
rect 35532 28704 35584 28756
rect 37280 28704 37332 28756
rect 37648 28704 37700 28756
rect 30564 28636 30616 28688
rect 32220 28636 32272 28688
rect 28724 28568 28776 28620
rect 31484 28568 31536 28620
rect 31852 28568 31904 28620
rect 25872 28500 25924 28552
rect 23480 28475 23532 28484
rect 18972 28364 19024 28416
rect 19984 28364 20036 28416
rect 23480 28441 23489 28475
rect 23489 28441 23523 28475
rect 23523 28441 23532 28475
rect 23480 28432 23532 28441
rect 23572 28432 23624 28484
rect 23940 28432 23992 28484
rect 26976 28500 27028 28552
rect 27160 28543 27212 28552
rect 27160 28509 27189 28543
rect 27189 28509 27212 28543
rect 27160 28500 27212 28509
rect 22008 28364 22060 28416
rect 23388 28364 23440 28416
rect 23756 28364 23808 28416
rect 24768 28364 24820 28416
rect 27068 28432 27120 28484
rect 28172 28543 28224 28552
rect 28172 28509 28181 28543
rect 28181 28509 28215 28543
rect 28215 28509 28224 28543
rect 28172 28500 28224 28509
rect 29460 28500 29512 28552
rect 30380 28500 30432 28552
rect 31024 28543 31076 28552
rect 31024 28509 31033 28543
rect 31033 28509 31067 28543
rect 31067 28509 31076 28543
rect 31024 28500 31076 28509
rect 32036 28500 32088 28552
rect 32220 28543 32272 28552
rect 32220 28509 32229 28543
rect 32229 28509 32263 28543
rect 32263 28509 32272 28543
rect 32220 28500 32272 28509
rect 33416 28568 33468 28620
rect 34336 28636 34388 28688
rect 34704 28636 34756 28688
rect 34796 28611 34848 28620
rect 34796 28577 34805 28611
rect 34805 28577 34839 28611
rect 34839 28577 34848 28611
rect 34796 28568 34848 28577
rect 33968 28543 34020 28552
rect 33968 28509 33977 28543
rect 33977 28509 34011 28543
rect 34011 28509 34020 28543
rect 33968 28500 34020 28509
rect 27252 28364 27304 28416
rect 28540 28432 28592 28484
rect 31852 28432 31904 28484
rect 32312 28432 32364 28484
rect 27988 28364 28040 28416
rect 30196 28364 30248 28416
rect 32220 28364 32272 28416
rect 32680 28364 32732 28416
rect 33876 28432 33928 28484
rect 34520 28500 34572 28552
rect 35900 28500 35952 28552
rect 36544 28500 36596 28552
rect 37280 28543 37332 28552
rect 37280 28509 37289 28543
rect 37289 28509 37323 28543
rect 37323 28509 37332 28543
rect 37280 28500 37332 28509
rect 35992 28475 36044 28484
rect 35992 28441 36001 28475
rect 36001 28441 36035 28475
rect 36035 28441 36044 28475
rect 35992 28432 36044 28441
rect 36544 28364 36596 28416
rect 37464 28432 37516 28484
rect 37924 28475 37976 28484
rect 37924 28441 37949 28475
rect 37949 28441 37976 28475
rect 37924 28432 37976 28441
rect 37372 28364 37424 28416
rect 38108 28407 38160 28416
rect 38108 28373 38117 28407
rect 38117 28373 38151 28407
rect 38151 28373 38160 28407
rect 38108 28364 38160 28373
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 16120 28160 16172 28212
rect 18236 28160 18288 28212
rect 17040 28092 17092 28144
rect 17132 28135 17184 28144
rect 17132 28101 17173 28135
rect 17173 28101 17184 28135
rect 17132 28092 17184 28101
rect 13820 28024 13872 28076
rect 14280 27956 14332 28008
rect 18328 28024 18380 28076
rect 19340 28092 19392 28144
rect 20628 28160 20680 28212
rect 24952 28160 25004 28212
rect 25044 28160 25096 28212
rect 25964 28160 26016 28212
rect 18972 28067 19024 28076
rect 18972 28033 18981 28067
rect 18981 28033 19015 28067
rect 19015 28033 19024 28067
rect 18972 28024 19024 28033
rect 19432 27999 19484 28008
rect 16856 27820 16908 27872
rect 17224 27820 17276 27872
rect 18696 27820 18748 27872
rect 19432 27965 19441 27999
rect 19441 27965 19475 27999
rect 19475 27965 19484 27999
rect 19432 27956 19484 27965
rect 19984 28024 20036 28076
rect 20628 28067 20680 28076
rect 20628 28033 20637 28067
rect 20637 28033 20671 28067
rect 20671 28033 20680 28067
rect 20628 28024 20680 28033
rect 20720 28067 20772 28076
rect 20720 28033 20729 28067
rect 20729 28033 20763 28067
rect 20763 28033 20772 28067
rect 20720 28024 20772 28033
rect 19708 27999 19760 28008
rect 19708 27965 19717 27999
rect 19717 27965 19751 27999
rect 19751 27965 19760 27999
rect 19708 27956 19760 27965
rect 20260 27956 20312 28008
rect 23020 28092 23072 28144
rect 28172 28160 28224 28212
rect 29552 28160 29604 28212
rect 30932 28160 30984 28212
rect 20996 28033 21005 28042
rect 21005 28033 21039 28042
rect 21039 28033 21048 28042
rect 20996 27990 21048 28033
rect 21180 28024 21232 28076
rect 22100 28024 22152 28076
rect 22744 28024 22796 28076
rect 24216 28024 24268 28076
rect 24768 28067 24820 28076
rect 24768 28033 24777 28067
rect 24777 28033 24811 28067
rect 24811 28033 24820 28067
rect 24768 28024 24820 28033
rect 25044 28024 25096 28076
rect 25228 28024 25280 28076
rect 28724 28092 28776 28144
rect 28816 28092 28868 28144
rect 31116 28135 31168 28144
rect 21272 27956 21324 28008
rect 23756 27956 23808 28008
rect 27712 28024 27764 28076
rect 28172 28024 28224 28076
rect 28908 28024 28960 28076
rect 31116 28101 31125 28135
rect 31125 28101 31159 28135
rect 31159 28101 31168 28135
rect 31116 28092 31168 28101
rect 31484 28160 31536 28212
rect 31852 28092 31904 28144
rect 32404 28135 32456 28144
rect 29184 28024 29236 28076
rect 28080 27956 28132 28008
rect 29368 28067 29420 28076
rect 29368 28033 29377 28067
rect 29377 28033 29411 28067
rect 29411 28033 29420 28067
rect 29368 28024 29420 28033
rect 29736 28024 29788 28076
rect 30840 28067 30892 28076
rect 29644 27956 29696 28008
rect 30840 28033 30849 28067
rect 30849 28033 30883 28067
rect 30883 28033 30892 28067
rect 30840 28024 30892 28033
rect 30932 28024 30984 28076
rect 31944 28024 31996 28076
rect 32404 28101 32413 28135
rect 32413 28101 32447 28135
rect 32447 28101 32456 28135
rect 32404 28092 32456 28101
rect 22376 27888 22428 27940
rect 26608 27888 26660 27940
rect 27620 27931 27672 27940
rect 27620 27897 27629 27931
rect 27629 27897 27663 27931
rect 27663 27897 27672 27931
rect 30104 27999 30156 28008
rect 30104 27965 30113 27999
rect 30113 27965 30147 27999
rect 30147 27965 30156 27999
rect 30104 27956 30156 27965
rect 30288 27956 30340 28008
rect 31392 27956 31444 28008
rect 27620 27888 27672 27897
rect 21824 27820 21876 27872
rect 22284 27820 22336 27872
rect 25780 27820 25832 27872
rect 25964 27820 26016 27872
rect 27436 27820 27488 27872
rect 28448 27820 28500 27872
rect 29000 27820 29052 27872
rect 29644 27820 29696 27872
rect 32036 27888 32088 27940
rect 32404 27888 32456 27940
rect 32772 28024 32824 28076
rect 32680 27888 32732 27940
rect 33600 28092 33652 28144
rect 33692 28067 33744 28076
rect 33692 28033 33701 28067
rect 33701 28033 33735 28067
rect 33735 28033 33744 28067
rect 33692 28024 33744 28033
rect 34428 28203 34480 28212
rect 34428 28169 34437 28203
rect 34437 28169 34471 28203
rect 34471 28169 34480 28203
rect 37648 28203 37700 28212
rect 34428 28160 34480 28169
rect 37648 28169 37657 28203
rect 37657 28169 37691 28203
rect 37691 28169 37700 28203
rect 37648 28160 37700 28169
rect 34520 28067 34572 28076
rect 34520 28033 34529 28067
rect 34529 28033 34563 28067
rect 34563 28033 34572 28067
rect 34520 28024 34572 28033
rect 33968 27956 34020 28008
rect 35440 28024 35492 28076
rect 35900 28067 35952 28076
rect 35900 28033 35909 28067
rect 35909 28033 35943 28067
rect 35943 28033 35952 28067
rect 35900 28024 35952 28033
rect 35992 28024 36044 28076
rect 36544 28067 36596 28076
rect 36544 28033 36553 28067
rect 36553 28033 36587 28067
rect 36587 28033 36596 28067
rect 36544 28024 36596 28033
rect 36636 27956 36688 28008
rect 37280 28024 37332 28076
rect 37464 28067 37516 28076
rect 37464 28033 37473 28067
rect 37473 28033 37507 28067
rect 37507 28033 37516 28067
rect 37464 28024 37516 28033
rect 37924 28024 37976 28076
rect 31944 27820 31996 27872
rect 33048 27820 33100 27872
rect 33876 27820 33928 27872
rect 36636 27863 36688 27872
rect 36636 27829 36645 27863
rect 36645 27829 36679 27863
rect 36679 27829 36688 27863
rect 36636 27820 36688 27829
rect 37740 27820 37792 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 16948 27659 17000 27668
rect 16948 27625 16957 27659
rect 16957 27625 16991 27659
rect 16991 27625 17000 27659
rect 16948 27616 17000 27625
rect 17776 27548 17828 27600
rect 19708 27616 19760 27668
rect 20352 27616 20404 27668
rect 20996 27616 21048 27668
rect 23020 27616 23072 27668
rect 25872 27659 25924 27668
rect 25872 27625 25881 27659
rect 25881 27625 25915 27659
rect 25915 27625 25924 27659
rect 25872 27616 25924 27625
rect 27896 27616 27948 27668
rect 20168 27548 20220 27600
rect 14280 27412 14332 27464
rect 14740 27455 14792 27464
rect 14740 27421 14749 27455
rect 14749 27421 14783 27455
rect 14783 27421 14792 27455
rect 14740 27412 14792 27421
rect 15936 27412 15988 27464
rect 17132 27480 17184 27532
rect 17224 27455 17276 27464
rect 17224 27421 17233 27455
rect 17233 27421 17267 27455
rect 17267 27421 17276 27455
rect 17224 27412 17276 27421
rect 18604 27480 18656 27532
rect 19340 27480 19392 27532
rect 18052 27455 18104 27464
rect 18052 27421 18061 27455
rect 18061 27421 18095 27455
rect 18095 27421 18104 27455
rect 18052 27412 18104 27421
rect 20168 27455 20220 27464
rect 16764 27344 16816 27396
rect 16856 27344 16908 27396
rect 19248 27344 19300 27396
rect 20168 27421 20177 27455
rect 20177 27421 20211 27455
rect 20211 27421 20220 27455
rect 20168 27412 20220 27421
rect 20628 27480 20680 27532
rect 24768 27548 24820 27600
rect 28080 27548 28132 27600
rect 28172 27548 28224 27600
rect 28448 27616 28500 27668
rect 31944 27616 31996 27668
rect 28540 27548 28592 27600
rect 28724 27548 28776 27600
rect 25504 27480 25556 27532
rect 20628 27344 20680 27396
rect 21088 27387 21140 27396
rect 21088 27353 21097 27387
rect 21097 27353 21131 27387
rect 21131 27353 21140 27387
rect 21088 27344 21140 27353
rect 21732 27344 21784 27396
rect 21916 27412 21968 27464
rect 23204 27455 23256 27464
rect 23204 27421 23213 27455
rect 23213 27421 23247 27455
rect 23247 27421 23256 27455
rect 23204 27412 23256 27421
rect 23940 27412 23992 27464
rect 24400 27412 24452 27464
rect 24952 27412 25004 27464
rect 26516 27455 26568 27464
rect 23020 27344 23072 27396
rect 23756 27344 23808 27396
rect 26516 27421 26525 27455
rect 26525 27421 26559 27455
rect 26559 27421 26568 27455
rect 26516 27412 26568 27421
rect 26700 27480 26752 27532
rect 31116 27548 31168 27600
rect 30748 27480 30800 27532
rect 31024 27480 31076 27532
rect 16120 27276 16172 27328
rect 17040 27276 17092 27328
rect 18512 27276 18564 27328
rect 20168 27276 20220 27328
rect 20536 27276 20588 27328
rect 22560 27276 22612 27328
rect 23296 27276 23348 27328
rect 24216 27276 24268 27328
rect 25688 27276 25740 27328
rect 26608 27319 26660 27328
rect 26608 27285 26617 27319
rect 26617 27285 26651 27319
rect 26651 27285 26660 27319
rect 26608 27276 26660 27285
rect 26884 27344 26936 27396
rect 27436 27412 27488 27464
rect 29368 27412 29420 27464
rect 29644 27455 29696 27464
rect 29644 27421 29653 27455
rect 29653 27421 29687 27455
rect 29687 27421 29696 27455
rect 29644 27412 29696 27421
rect 29736 27412 29788 27464
rect 30380 27412 30432 27464
rect 30472 27455 30524 27464
rect 30472 27421 30481 27455
rect 30481 27421 30515 27455
rect 30515 27421 30524 27455
rect 30472 27412 30524 27421
rect 30656 27412 30708 27464
rect 30840 27412 30892 27464
rect 27712 27387 27764 27396
rect 27712 27353 27721 27387
rect 27721 27353 27755 27387
rect 27755 27353 27764 27387
rect 27712 27344 27764 27353
rect 27988 27344 28040 27396
rect 31852 27548 31904 27600
rect 32312 27574 32364 27626
rect 32404 27574 32456 27626
rect 32496 27616 32548 27668
rect 34520 27616 34572 27668
rect 28356 27319 28408 27328
rect 28356 27285 28381 27319
rect 28381 27285 28408 27319
rect 28356 27276 28408 27285
rect 28540 27319 28592 27328
rect 28540 27285 28549 27319
rect 28549 27285 28583 27319
rect 28583 27285 28592 27319
rect 30380 27319 30432 27328
rect 28540 27276 28592 27285
rect 30380 27285 30389 27319
rect 30389 27285 30423 27319
rect 30423 27285 30432 27319
rect 30380 27276 30432 27285
rect 30472 27276 30524 27328
rect 31944 27480 31996 27532
rect 32036 27480 32088 27532
rect 31484 27412 31536 27464
rect 31852 27412 31904 27464
rect 37464 27548 37516 27600
rect 34428 27480 34480 27532
rect 31760 27344 31812 27396
rect 33232 27412 33284 27464
rect 34612 27412 34664 27464
rect 35992 27480 36044 27532
rect 36176 27523 36228 27532
rect 36176 27489 36185 27523
rect 36185 27489 36219 27523
rect 36219 27489 36228 27523
rect 36176 27480 36228 27489
rect 36728 27480 36780 27532
rect 35624 27455 35676 27464
rect 35624 27421 35633 27455
rect 35633 27421 35667 27455
rect 35667 27421 35676 27455
rect 35624 27412 35676 27421
rect 36360 27412 36412 27464
rect 37740 27455 37792 27464
rect 37740 27421 37749 27455
rect 37749 27421 37783 27455
rect 37783 27421 37792 27455
rect 37740 27412 37792 27421
rect 38108 27412 38160 27464
rect 31484 27276 31536 27328
rect 33416 27276 33468 27328
rect 33692 27319 33744 27328
rect 33692 27285 33701 27319
rect 33701 27285 33735 27319
rect 33735 27285 33744 27319
rect 33692 27276 33744 27285
rect 33784 27276 33836 27328
rect 35072 27276 35124 27328
rect 36084 27276 36136 27328
rect 37280 27276 37332 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 15936 27072 15988 27124
rect 20260 27072 20312 27124
rect 20352 27115 20404 27124
rect 20352 27081 20361 27115
rect 20361 27081 20395 27115
rect 20395 27081 20404 27115
rect 20352 27072 20404 27081
rect 24860 27072 24912 27124
rect 25228 27072 25280 27124
rect 26056 27072 26108 27124
rect 18052 27047 18104 27056
rect 18052 27013 18061 27047
rect 18061 27013 18095 27047
rect 18095 27013 18104 27047
rect 18052 27004 18104 27013
rect 20996 27004 21048 27056
rect 22008 27004 22060 27056
rect 14648 26979 14700 26988
rect 14648 26945 14657 26979
rect 14657 26945 14691 26979
rect 14691 26945 14700 26979
rect 14648 26936 14700 26945
rect 15936 26979 15988 26988
rect 15936 26945 15945 26979
rect 15945 26945 15979 26979
rect 15979 26945 15988 26979
rect 15936 26936 15988 26945
rect 16120 26979 16172 26988
rect 16120 26945 16129 26979
rect 16129 26945 16163 26979
rect 16163 26945 16172 26979
rect 16120 26936 16172 26945
rect 16764 26979 16816 26988
rect 16764 26945 16773 26979
rect 16773 26945 16807 26979
rect 16807 26945 16816 26979
rect 16764 26936 16816 26945
rect 17960 26936 18012 26988
rect 19248 26936 19300 26988
rect 14280 26868 14332 26920
rect 15292 26868 15344 26920
rect 19524 26868 19576 26920
rect 18144 26800 18196 26852
rect 18328 26800 18380 26852
rect 20076 26936 20128 26988
rect 20444 26979 20496 26988
rect 20444 26945 20453 26979
rect 20453 26945 20487 26979
rect 20487 26945 20496 26979
rect 20444 26936 20496 26945
rect 20628 26936 20680 26988
rect 22376 26979 22428 26988
rect 22376 26945 22385 26979
rect 22385 26945 22419 26979
rect 22419 26945 22428 26979
rect 22376 26936 22428 26945
rect 24676 27004 24728 27056
rect 25412 27004 25464 27056
rect 28448 27047 28500 27056
rect 28448 27013 28457 27047
rect 28457 27013 28491 27047
rect 28491 27013 28500 27047
rect 28448 27004 28500 27013
rect 33048 27072 33100 27124
rect 33140 27072 33192 27124
rect 29736 27004 29788 27056
rect 30104 27004 30156 27056
rect 32496 27047 32548 27056
rect 32496 27013 32505 27047
rect 32505 27013 32539 27047
rect 32539 27013 32548 27047
rect 32496 27004 32548 27013
rect 33324 27004 33376 27056
rect 33692 27004 33744 27056
rect 33876 27072 33928 27124
rect 23572 26936 23624 26988
rect 23756 26936 23808 26988
rect 24584 26936 24636 26988
rect 24952 26979 25004 26988
rect 24952 26945 24961 26979
rect 24961 26945 24995 26979
rect 24995 26945 25004 26979
rect 24952 26936 25004 26945
rect 25320 26936 25372 26988
rect 25504 26936 25556 26988
rect 25780 26979 25832 26988
rect 25780 26945 25789 26979
rect 25789 26945 25823 26979
rect 25823 26945 25832 26979
rect 25780 26936 25832 26945
rect 27528 26936 27580 26988
rect 28080 26936 28132 26988
rect 29644 26979 29696 26988
rect 20260 26868 20312 26920
rect 22744 26911 22796 26920
rect 22744 26877 22753 26911
rect 22753 26877 22787 26911
rect 22787 26877 22796 26911
rect 22744 26868 22796 26877
rect 23020 26868 23072 26920
rect 25688 26868 25740 26920
rect 19984 26800 20036 26852
rect 25412 26800 25464 26852
rect 26976 26911 27028 26920
rect 26976 26877 26985 26911
rect 26985 26877 27019 26911
rect 27019 26877 27028 26911
rect 26976 26868 27028 26877
rect 27436 26868 27488 26920
rect 28356 26868 28408 26920
rect 29644 26945 29653 26979
rect 29653 26945 29687 26979
rect 29687 26945 29696 26979
rect 29644 26936 29696 26945
rect 30012 26979 30064 26988
rect 28816 26868 28868 26920
rect 29000 26868 29052 26920
rect 29460 26868 29512 26920
rect 30012 26945 30021 26979
rect 30021 26945 30055 26979
rect 30055 26945 30064 26979
rect 30012 26936 30064 26945
rect 30564 26936 30616 26988
rect 30656 26911 30708 26920
rect 30656 26877 30665 26911
rect 30665 26877 30699 26911
rect 30699 26877 30708 26911
rect 30656 26868 30708 26877
rect 30840 26936 30892 26988
rect 32220 26936 32272 26988
rect 31392 26868 31444 26920
rect 31576 26868 31628 26920
rect 31760 26868 31812 26920
rect 32404 26979 32456 26988
rect 32404 26945 32413 26979
rect 32413 26945 32447 26979
rect 32447 26945 32456 26979
rect 32404 26936 32456 26945
rect 34612 26979 34664 26988
rect 34612 26945 34621 26979
rect 34621 26945 34655 26979
rect 34655 26945 34664 26979
rect 34612 26936 34664 26945
rect 35624 27004 35676 27056
rect 33508 26868 33560 26920
rect 31852 26800 31904 26852
rect 33048 26800 33100 26852
rect 34428 26868 34480 26920
rect 16672 26732 16724 26784
rect 16856 26775 16908 26784
rect 16856 26741 16865 26775
rect 16865 26741 16899 26775
rect 16899 26741 16908 26775
rect 16856 26732 16908 26741
rect 17592 26732 17644 26784
rect 17776 26732 17828 26784
rect 17960 26732 18012 26784
rect 18236 26775 18288 26784
rect 18236 26741 18245 26775
rect 18245 26741 18279 26775
rect 18279 26741 18288 26775
rect 18236 26732 18288 26741
rect 19892 26732 19944 26784
rect 24308 26732 24360 26784
rect 27528 26732 27580 26784
rect 28448 26732 28500 26784
rect 29092 26732 29144 26784
rect 30564 26732 30616 26784
rect 31484 26732 31536 26784
rect 33232 26732 33284 26784
rect 34520 26800 34572 26852
rect 35072 26936 35124 26988
rect 35716 26979 35768 26988
rect 35716 26945 35725 26979
rect 35725 26945 35759 26979
rect 35759 26945 35768 26979
rect 35716 26936 35768 26945
rect 35900 26979 35952 26988
rect 35900 26945 35909 26979
rect 35909 26945 35943 26979
rect 35943 26945 35952 26979
rect 36452 26979 36504 26988
rect 35900 26936 35952 26945
rect 36452 26945 36461 26979
rect 36461 26945 36495 26979
rect 36495 26945 36504 26979
rect 36452 26936 36504 26945
rect 36544 26936 36596 26988
rect 37188 26936 37240 26988
rect 35624 26911 35676 26920
rect 35624 26877 35633 26911
rect 35633 26877 35667 26911
rect 35667 26877 35676 26911
rect 35624 26868 35676 26877
rect 37372 26911 37424 26920
rect 37372 26877 37381 26911
rect 37381 26877 37415 26911
rect 37415 26877 37424 26911
rect 37372 26868 37424 26877
rect 36728 26800 36780 26852
rect 35348 26732 35400 26784
rect 36452 26732 36504 26784
rect 37740 26775 37792 26784
rect 37740 26741 37749 26775
rect 37749 26741 37783 26775
rect 37783 26741 37792 26775
rect 37740 26732 37792 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 14280 26528 14332 26580
rect 15476 26528 15528 26580
rect 16764 26571 16816 26580
rect 16764 26537 16773 26571
rect 16773 26537 16807 26571
rect 16807 26537 16816 26571
rect 16764 26528 16816 26537
rect 17776 26571 17828 26580
rect 17776 26537 17785 26571
rect 17785 26537 17819 26571
rect 17819 26537 17828 26571
rect 17776 26528 17828 26537
rect 14372 26324 14424 26376
rect 15292 26367 15344 26376
rect 15292 26333 15301 26367
rect 15301 26333 15335 26367
rect 15335 26333 15344 26367
rect 15292 26324 15344 26333
rect 15476 26324 15528 26376
rect 14004 26256 14056 26308
rect 16672 26324 16724 26376
rect 18236 26392 18288 26444
rect 19340 26460 19392 26512
rect 21272 26392 21324 26444
rect 21456 26435 21508 26444
rect 21456 26401 21465 26435
rect 21465 26401 21499 26435
rect 21499 26401 21508 26435
rect 21456 26392 21508 26401
rect 21916 26528 21968 26580
rect 24124 26528 24176 26580
rect 26884 26528 26936 26580
rect 27712 26528 27764 26580
rect 27804 26528 27856 26580
rect 22468 26460 22520 26512
rect 25320 26460 25372 26512
rect 26424 26460 26476 26512
rect 28172 26460 28224 26512
rect 31760 26528 31812 26580
rect 33416 26528 33468 26580
rect 35900 26571 35952 26580
rect 30656 26460 30708 26512
rect 31576 26460 31628 26512
rect 24216 26392 24268 26444
rect 19892 26367 19944 26376
rect 16120 26256 16172 26308
rect 19892 26333 19901 26367
rect 19901 26333 19935 26367
rect 19935 26333 19944 26367
rect 19892 26324 19944 26333
rect 20168 26367 20220 26376
rect 20168 26333 20177 26367
rect 20177 26333 20211 26367
rect 20211 26333 20220 26367
rect 20168 26324 20220 26333
rect 20720 26324 20772 26376
rect 20996 26324 21048 26376
rect 21916 26367 21968 26376
rect 21916 26333 21925 26367
rect 21925 26333 21959 26367
rect 21959 26333 21968 26367
rect 21916 26324 21968 26333
rect 23388 26324 23440 26376
rect 24308 26324 24360 26376
rect 20076 26256 20128 26308
rect 24400 26256 24452 26308
rect 27068 26324 27120 26376
rect 29000 26392 29052 26444
rect 29184 26392 29236 26444
rect 27528 26367 27580 26376
rect 27528 26333 27537 26367
rect 27537 26333 27571 26367
rect 27571 26333 27580 26367
rect 27528 26324 27580 26333
rect 27804 26367 27856 26376
rect 27804 26333 27813 26367
rect 27813 26333 27847 26367
rect 27847 26333 27856 26367
rect 27804 26324 27856 26333
rect 28540 26324 28592 26376
rect 30012 26324 30064 26376
rect 30472 26367 30524 26376
rect 30472 26333 30481 26367
rect 30481 26333 30515 26367
rect 30515 26333 30524 26367
rect 30472 26324 30524 26333
rect 30656 26324 30708 26376
rect 28816 26256 28868 26308
rect 29000 26256 29052 26308
rect 30380 26256 30432 26308
rect 31024 26392 31076 26444
rect 31944 26392 31996 26444
rect 32588 26392 32640 26444
rect 34336 26460 34388 26512
rect 34520 26460 34572 26512
rect 34980 26460 35032 26512
rect 35900 26537 35909 26571
rect 35909 26537 35943 26571
rect 35943 26537 35952 26571
rect 35900 26528 35952 26537
rect 36176 26571 36228 26580
rect 36176 26537 36185 26571
rect 36185 26537 36219 26571
rect 36219 26537 36228 26571
rect 36176 26528 36228 26537
rect 37556 26460 37608 26512
rect 32496 26367 32548 26376
rect 32496 26333 32505 26367
rect 32505 26333 32539 26367
rect 32539 26333 32548 26367
rect 32496 26324 32548 26333
rect 32772 26367 32824 26376
rect 31852 26299 31904 26308
rect 31852 26265 31861 26299
rect 31861 26265 31895 26299
rect 31895 26265 31904 26299
rect 32772 26333 32781 26367
rect 32781 26333 32815 26367
rect 32815 26333 32824 26367
rect 32772 26324 32824 26333
rect 33876 26392 33928 26444
rect 34060 26392 34112 26444
rect 35624 26392 35676 26444
rect 33508 26324 33560 26376
rect 34796 26324 34848 26376
rect 34980 26367 35032 26376
rect 34980 26333 34989 26367
rect 34989 26333 35023 26367
rect 35023 26333 35032 26367
rect 34980 26324 35032 26333
rect 31852 26256 31904 26265
rect 21364 26188 21416 26240
rect 21732 26231 21784 26240
rect 21732 26197 21741 26231
rect 21741 26197 21775 26231
rect 21775 26197 21784 26231
rect 21732 26188 21784 26197
rect 23020 26188 23072 26240
rect 27252 26188 27304 26240
rect 33232 26256 33284 26308
rect 34612 26256 34664 26308
rect 35532 26324 35584 26376
rect 36452 26324 36504 26376
rect 37740 26367 37792 26376
rect 37740 26333 37749 26367
rect 37749 26333 37783 26367
rect 37783 26333 37792 26367
rect 37740 26324 37792 26333
rect 37372 26256 37424 26308
rect 33048 26188 33100 26240
rect 33508 26188 33560 26240
rect 36544 26188 36596 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 14372 25984 14424 26036
rect 14648 25984 14700 26036
rect 16120 26027 16172 26036
rect 16120 25993 16129 26027
rect 16129 25993 16163 26027
rect 16163 25993 16172 26027
rect 16120 25984 16172 25993
rect 17960 25984 18012 26036
rect 18512 25984 18564 26036
rect 21456 25984 21508 26036
rect 25596 25984 25648 26036
rect 25872 25984 25924 26036
rect 26608 25984 26660 26036
rect 28356 25984 28408 26036
rect 30012 25984 30064 26036
rect 13912 25848 13964 25900
rect 15200 25916 15252 25968
rect 18144 25916 18196 25968
rect 14648 25891 14700 25900
rect 14648 25857 14657 25891
rect 14657 25857 14691 25891
rect 14691 25857 14700 25891
rect 14648 25848 14700 25857
rect 15384 25891 15436 25900
rect 15384 25857 15393 25891
rect 15393 25857 15427 25891
rect 15427 25857 15436 25891
rect 15384 25848 15436 25857
rect 15752 25848 15804 25900
rect 19248 25916 19300 25968
rect 20076 25848 20128 25900
rect 20168 25848 20220 25900
rect 25504 25916 25556 25968
rect 27436 25959 27488 25968
rect 21364 25848 21416 25900
rect 22376 25891 22428 25900
rect 22376 25857 22385 25891
rect 22385 25857 22419 25891
rect 22419 25857 22428 25891
rect 22376 25848 22428 25857
rect 23020 25848 23072 25900
rect 23940 25848 23992 25900
rect 13820 25755 13872 25764
rect 13820 25721 13829 25755
rect 13829 25721 13863 25755
rect 13863 25721 13872 25755
rect 13820 25712 13872 25721
rect 16396 25780 16448 25832
rect 19984 25780 20036 25832
rect 21916 25780 21968 25832
rect 22284 25780 22336 25832
rect 24584 25848 24636 25900
rect 24400 25780 24452 25832
rect 20352 25712 20404 25764
rect 23388 25712 23440 25764
rect 23848 25712 23900 25764
rect 25228 25780 25280 25832
rect 25872 25891 25924 25900
rect 25872 25857 25881 25891
rect 25881 25857 25915 25891
rect 25915 25857 25924 25891
rect 25872 25848 25924 25857
rect 26056 25848 26108 25900
rect 27436 25925 27445 25959
rect 27445 25925 27479 25959
rect 27479 25925 27488 25959
rect 27436 25916 27488 25925
rect 27988 25916 28040 25968
rect 28908 25916 28960 25968
rect 29092 25916 29144 25968
rect 29368 25959 29420 25968
rect 29368 25925 29377 25959
rect 29377 25925 29411 25959
rect 29411 25925 29420 25959
rect 29368 25916 29420 25925
rect 26516 25848 26568 25900
rect 26792 25848 26844 25900
rect 29736 25848 29788 25900
rect 30104 25848 30156 25900
rect 30288 25848 30340 25900
rect 32036 25984 32088 26036
rect 32496 25984 32548 26036
rect 33784 25984 33836 26036
rect 36728 25984 36780 26036
rect 30932 25916 30984 25968
rect 30840 25848 30892 25900
rect 31024 25848 31076 25900
rect 31300 25891 31352 25900
rect 31300 25857 31309 25891
rect 31309 25857 31343 25891
rect 31343 25857 31352 25891
rect 31300 25848 31352 25857
rect 26240 25780 26292 25832
rect 28632 25780 28684 25832
rect 28816 25823 28868 25832
rect 28816 25789 28825 25823
rect 28825 25789 28859 25823
rect 28859 25789 28868 25823
rect 28816 25780 28868 25789
rect 31392 25780 31444 25832
rect 31944 25916 31996 25968
rect 32772 25916 32824 25968
rect 33508 25959 33560 25968
rect 33508 25925 33517 25959
rect 33517 25925 33551 25959
rect 33551 25925 33560 25959
rect 33508 25916 33560 25925
rect 35716 25916 35768 25968
rect 32312 25891 32364 25900
rect 32312 25857 32321 25891
rect 32321 25857 32355 25891
rect 32355 25857 32364 25891
rect 32312 25848 32364 25857
rect 32956 25848 33008 25900
rect 33140 25848 33192 25900
rect 34336 25891 34388 25900
rect 34336 25857 34345 25891
rect 34345 25857 34379 25891
rect 34379 25857 34388 25891
rect 34336 25848 34388 25857
rect 35992 25848 36044 25900
rect 36176 25891 36228 25900
rect 36176 25857 36185 25891
rect 36185 25857 36219 25891
rect 36219 25857 36228 25891
rect 36176 25848 36228 25857
rect 37464 25891 37516 25900
rect 37464 25857 37473 25891
rect 37473 25857 37507 25891
rect 37507 25857 37516 25891
rect 37464 25848 37516 25857
rect 37556 25823 37608 25832
rect 37556 25789 37565 25823
rect 37565 25789 37599 25823
rect 37599 25789 37608 25823
rect 37556 25780 37608 25789
rect 25872 25712 25924 25764
rect 26056 25755 26108 25764
rect 26056 25721 26065 25755
rect 26065 25721 26099 25755
rect 26099 25721 26108 25755
rect 26056 25712 26108 25721
rect 27804 25712 27856 25764
rect 30656 25712 30708 25764
rect 31668 25712 31720 25764
rect 15476 25644 15528 25696
rect 18328 25644 18380 25696
rect 19064 25687 19116 25696
rect 19064 25653 19073 25687
rect 19073 25653 19107 25687
rect 19107 25653 19116 25687
rect 19064 25644 19116 25653
rect 23112 25644 23164 25696
rect 23572 25644 23624 25696
rect 25596 25644 25648 25696
rect 26424 25644 26476 25696
rect 28540 25644 28592 25696
rect 29920 25644 29972 25696
rect 30288 25644 30340 25696
rect 30748 25644 30800 25696
rect 31392 25644 31444 25696
rect 32496 25644 32548 25696
rect 33876 25687 33928 25696
rect 33876 25653 33885 25687
rect 33885 25653 33919 25687
rect 33919 25653 33928 25687
rect 33876 25644 33928 25653
rect 34520 25687 34572 25696
rect 34520 25653 34529 25687
rect 34529 25653 34563 25687
rect 34563 25653 34572 25687
rect 34520 25644 34572 25653
rect 35900 25687 35952 25696
rect 35900 25653 35909 25687
rect 35909 25653 35943 25687
rect 35943 25653 35952 25687
rect 35900 25644 35952 25653
rect 37556 25644 37608 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 14004 25440 14056 25492
rect 14740 25440 14792 25492
rect 15384 25440 15436 25492
rect 15752 25483 15804 25492
rect 15752 25449 15761 25483
rect 15761 25449 15795 25483
rect 15795 25449 15804 25483
rect 15752 25440 15804 25449
rect 18052 25440 18104 25492
rect 21088 25440 21140 25492
rect 24768 25440 24820 25492
rect 24860 25440 24912 25492
rect 20720 25372 20772 25424
rect 22652 25372 22704 25424
rect 23388 25372 23440 25424
rect 23480 25372 23532 25424
rect 31024 25440 31076 25492
rect 31208 25440 31260 25492
rect 34796 25440 34848 25492
rect 36176 25440 36228 25492
rect 15384 25304 15436 25356
rect 16396 25347 16448 25356
rect 16396 25313 16405 25347
rect 16405 25313 16439 25347
rect 16439 25313 16448 25347
rect 16396 25304 16448 25313
rect 21916 25304 21968 25356
rect 22836 25347 22888 25356
rect 14096 25236 14148 25288
rect 14280 25279 14332 25288
rect 14280 25245 14289 25279
rect 14289 25245 14323 25279
rect 14323 25245 14332 25279
rect 14280 25236 14332 25245
rect 15292 25279 15344 25288
rect 15292 25245 15301 25279
rect 15301 25245 15335 25279
rect 15335 25245 15344 25279
rect 15292 25236 15344 25245
rect 16120 25236 16172 25288
rect 16672 25279 16724 25288
rect 16672 25245 16681 25279
rect 16681 25245 16715 25279
rect 16715 25245 16724 25279
rect 16672 25236 16724 25245
rect 17960 25236 18012 25288
rect 19432 25236 19484 25288
rect 20076 25236 20128 25288
rect 20996 25236 21048 25288
rect 22836 25313 22845 25347
rect 22845 25313 22879 25347
rect 22879 25313 22888 25347
rect 22836 25304 22888 25313
rect 23848 25347 23900 25356
rect 23848 25313 23857 25347
rect 23857 25313 23891 25347
rect 23891 25313 23900 25347
rect 23848 25304 23900 25313
rect 25872 25304 25924 25356
rect 27620 25304 27672 25356
rect 22560 25279 22612 25288
rect 22560 25245 22569 25279
rect 22569 25245 22603 25279
rect 22603 25245 22612 25279
rect 22560 25236 22612 25245
rect 21364 25168 21416 25220
rect 23756 25236 23808 25288
rect 24400 25279 24452 25288
rect 24400 25245 24409 25279
rect 24409 25245 24443 25279
rect 24443 25245 24452 25279
rect 24400 25236 24452 25245
rect 24676 25279 24728 25288
rect 24676 25245 24685 25279
rect 24685 25245 24719 25279
rect 24719 25245 24728 25279
rect 24676 25236 24728 25245
rect 24124 25168 24176 25220
rect 26516 25236 26568 25288
rect 26884 25279 26936 25288
rect 26884 25245 26893 25279
rect 26893 25245 26927 25279
rect 26927 25245 26936 25279
rect 26884 25236 26936 25245
rect 27068 25279 27120 25288
rect 27068 25245 27077 25279
rect 27077 25245 27111 25279
rect 27111 25245 27120 25279
rect 27068 25236 27120 25245
rect 26700 25168 26752 25220
rect 28816 25372 28868 25424
rect 30380 25372 30432 25424
rect 28080 25236 28132 25288
rect 28632 25304 28684 25356
rect 30012 25304 30064 25356
rect 28540 25279 28592 25288
rect 28540 25245 28549 25279
rect 28549 25245 28583 25279
rect 28583 25245 28592 25279
rect 28540 25236 28592 25245
rect 29460 25236 29512 25288
rect 29092 25168 29144 25220
rect 30656 25236 30708 25288
rect 31208 25236 31260 25288
rect 31300 25168 31352 25220
rect 34060 25304 34112 25356
rect 34520 25304 34572 25356
rect 37556 25347 37608 25356
rect 37556 25313 37565 25347
rect 37565 25313 37599 25347
rect 37599 25313 37608 25347
rect 37556 25304 37608 25313
rect 32312 25236 32364 25288
rect 32864 25236 32916 25288
rect 35256 25279 35308 25288
rect 35256 25245 35265 25279
rect 35265 25245 35299 25279
rect 35299 25245 35308 25279
rect 35256 25236 35308 25245
rect 37832 25236 37884 25288
rect 18604 25100 18656 25152
rect 23388 25100 23440 25152
rect 23572 25100 23624 25152
rect 25872 25143 25924 25152
rect 25872 25109 25881 25143
rect 25881 25109 25915 25143
rect 25915 25109 25924 25143
rect 25872 25100 25924 25109
rect 26516 25100 26568 25152
rect 27620 25100 27672 25152
rect 30656 25100 30708 25152
rect 30748 25143 30800 25152
rect 30748 25109 30773 25143
rect 30773 25109 30800 25143
rect 30932 25143 30984 25152
rect 30748 25100 30800 25109
rect 30932 25109 30941 25143
rect 30941 25109 30975 25143
rect 30975 25109 30984 25143
rect 30932 25100 30984 25109
rect 35716 25168 35768 25220
rect 32220 25100 32272 25152
rect 33692 25100 33744 25152
rect 35992 25143 36044 25152
rect 35992 25109 36017 25143
rect 36017 25109 36044 25143
rect 36176 25143 36228 25152
rect 35992 25100 36044 25109
rect 36176 25109 36185 25143
rect 36185 25109 36219 25143
rect 36219 25109 36228 25143
rect 36176 25100 36228 25109
rect 37556 25100 37608 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 14280 24896 14332 24948
rect 18972 24896 19024 24948
rect 19064 24896 19116 24948
rect 24308 24896 24360 24948
rect 24400 24896 24452 24948
rect 26240 24896 26292 24948
rect 31576 24896 31628 24948
rect 31944 24896 31996 24948
rect 34060 24939 34112 24948
rect 34060 24905 34069 24939
rect 34069 24905 34103 24939
rect 34103 24905 34112 24939
rect 34060 24896 34112 24905
rect 37464 24896 37516 24948
rect 12992 24828 13044 24880
rect 13820 24828 13872 24880
rect 15016 24871 15068 24880
rect 14280 24760 14332 24812
rect 15016 24837 15025 24871
rect 15025 24837 15059 24871
rect 15059 24837 15068 24871
rect 15016 24828 15068 24837
rect 10048 24692 10100 24744
rect 15016 24692 15068 24744
rect 15200 24692 15252 24744
rect 15936 24760 15988 24812
rect 18052 24760 18104 24812
rect 18604 24803 18656 24812
rect 18604 24769 18613 24803
rect 18613 24769 18647 24803
rect 18647 24769 18656 24803
rect 18604 24760 18656 24769
rect 19800 24760 19852 24812
rect 20444 24803 20496 24812
rect 20444 24769 20453 24803
rect 20453 24769 20487 24803
rect 20487 24769 20496 24803
rect 20444 24760 20496 24769
rect 20536 24803 20588 24812
rect 20536 24769 20545 24803
rect 20545 24769 20579 24803
rect 20579 24769 20588 24803
rect 20536 24760 20588 24769
rect 21180 24760 21232 24812
rect 21272 24803 21324 24812
rect 21272 24769 21281 24803
rect 21281 24769 21315 24803
rect 21315 24769 21324 24803
rect 21272 24760 21324 24769
rect 14648 24624 14700 24676
rect 16764 24692 16816 24744
rect 21732 24760 21784 24812
rect 23020 24760 23072 24812
rect 24676 24828 24728 24880
rect 25228 24828 25280 24880
rect 26056 24828 26108 24880
rect 23848 24760 23900 24812
rect 25504 24760 25556 24812
rect 25964 24760 26016 24812
rect 26240 24760 26292 24812
rect 26792 24760 26844 24812
rect 27528 24828 27580 24880
rect 28264 24828 28316 24880
rect 28080 24803 28132 24812
rect 16672 24624 16724 24676
rect 15200 24599 15252 24608
rect 15200 24565 15209 24599
rect 15209 24565 15243 24599
rect 15243 24565 15252 24599
rect 15200 24556 15252 24565
rect 18144 24624 18196 24676
rect 17776 24556 17828 24608
rect 19432 24624 19484 24676
rect 22560 24692 22612 24744
rect 24860 24692 24912 24744
rect 25872 24692 25924 24744
rect 26424 24735 26476 24744
rect 26424 24701 26433 24735
rect 26433 24701 26467 24735
rect 26467 24701 26476 24735
rect 26424 24692 26476 24701
rect 28080 24769 28089 24803
rect 28089 24769 28123 24803
rect 28123 24769 28132 24803
rect 28080 24760 28132 24769
rect 28908 24803 28960 24812
rect 28908 24769 28917 24803
rect 28917 24769 28951 24803
rect 28951 24769 28960 24803
rect 31024 24828 31076 24880
rect 31300 24828 31352 24880
rect 28908 24760 28960 24769
rect 27252 24692 27304 24744
rect 30380 24735 30432 24744
rect 30380 24701 30389 24735
rect 30389 24701 30423 24735
rect 30423 24701 30432 24735
rect 30380 24692 30432 24701
rect 30656 24760 30708 24812
rect 31208 24735 31260 24744
rect 31208 24701 31217 24735
rect 31217 24701 31251 24735
rect 31251 24701 31260 24735
rect 31208 24692 31260 24701
rect 32036 24760 32088 24812
rect 33140 24828 33192 24880
rect 35256 24828 35308 24880
rect 35900 24871 35952 24880
rect 35900 24837 35909 24871
rect 35909 24837 35943 24871
rect 35943 24837 35952 24871
rect 35900 24828 35952 24837
rect 32772 24803 32824 24812
rect 32772 24769 32781 24803
rect 32781 24769 32815 24803
rect 32815 24769 32824 24803
rect 32772 24760 32824 24769
rect 33876 24760 33928 24812
rect 34336 24760 34388 24812
rect 21272 24624 21324 24676
rect 23480 24667 23532 24676
rect 20720 24556 20772 24608
rect 21824 24556 21876 24608
rect 23480 24633 23489 24667
rect 23489 24633 23523 24667
rect 23523 24633 23532 24667
rect 23480 24624 23532 24633
rect 29276 24667 29328 24676
rect 29276 24633 29285 24667
rect 29285 24633 29319 24667
rect 29319 24633 29328 24667
rect 29276 24624 29328 24633
rect 32036 24624 32088 24676
rect 33784 24692 33836 24744
rect 35992 24760 36044 24812
rect 36728 24760 36780 24812
rect 36176 24692 36228 24744
rect 37188 24692 37240 24744
rect 37740 24803 37792 24812
rect 37740 24769 37749 24803
rect 37749 24769 37783 24803
rect 37783 24769 37792 24803
rect 37740 24760 37792 24769
rect 32772 24624 32824 24676
rect 34796 24624 34848 24676
rect 22744 24556 22796 24608
rect 23112 24556 23164 24608
rect 23664 24556 23716 24608
rect 23756 24556 23808 24608
rect 26240 24599 26292 24608
rect 26240 24565 26249 24599
rect 26249 24565 26283 24599
rect 26283 24565 26292 24599
rect 26240 24556 26292 24565
rect 26792 24556 26844 24608
rect 27068 24556 27120 24608
rect 31576 24556 31628 24608
rect 31852 24556 31904 24608
rect 32404 24556 32456 24608
rect 35440 24556 35492 24608
rect 36268 24599 36320 24608
rect 36268 24565 36277 24599
rect 36277 24565 36311 24599
rect 36311 24565 36320 24599
rect 36268 24556 36320 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 13912 24284 13964 24336
rect 16120 24395 16172 24404
rect 15200 24284 15252 24336
rect 15292 24327 15344 24336
rect 15292 24293 15301 24327
rect 15301 24293 15335 24327
rect 15335 24293 15344 24327
rect 16120 24361 16129 24395
rect 16129 24361 16163 24395
rect 16163 24361 16172 24395
rect 16120 24352 16172 24361
rect 16488 24352 16540 24404
rect 19432 24352 19484 24404
rect 19800 24395 19852 24404
rect 19800 24361 19809 24395
rect 19809 24361 19843 24395
rect 19843 24361 19852 24395
rect 19800 24352 19852 24361
rect 20444 24352 20496 24404
rect 15292 24284 15344 24293
rect 10232 24216 10284 24268
rect 14096 24216 14148 24268
rect 20168 24216 20220 24268
rect 20444 24216 20496 24268
rect 11612 24191 11664 24200
rect 11612 24157 11621 24191
rect 11621 24157 11655 24191
rect 11655 24157 11664 24191
rect 11612 24148 11664 24157
rect 11888 24148 11940 24200
rect 17500 24191 17552 24200
rect 10324 24080 10376 24132
rect 17500 24157 17509 24191
rect 17509 24157 17543 24191
rect 17543 24157 17552 24191
rect 17500 24148 17552 24157
rect 18512 24191 18564 24200
rect 14280 24123 14332 24132
rect 14280 24089 14310 24123
rect 14310 24089 14332 24123
rect 14280 24080 14332 24089
rect 15016 24080 15068 24132
rect 15660 24080 15712 24132
rect 15844 24080 15896 24132
rect 16764 24123 16816 24132
rect 16764 24089 16789 24123
rect 16789 24089 16816 24123
rect 16764 24080 16816 24089
rect 13452 24012 13504 24064
rect 14464 24012 14516 24064
rect 15108 24055 15160 24064
rect 15108 24021 15133 24055
rect 15133 24021 15160 24055
rect 15108 24012 15160 24021
rect 18236 24012 18288 24064
rect 18512 24157 18521 24191
rect 18521 24157 18555 24191
rect 18555 24157 18564 24191
rect 18512 24148 18564 24157
rect 22192 24352 22244 24404
rect 26240 24352 26292 24404
rect 26884 24352 26936 24404
rect 27436 24284 27488 24336
rect 22376 24216 22428 24268
rect 23480 24216 23532 24268
rect 24124 24216 24176 24268
rect 20996 24191 21048 24200
rect 20444 24123 20496 24132
rect 20444 24089 20453 24123
rect 20453 24089 20487 24123
rect 20487 24089 20496 24123
rect 20444 24080 20496 24089
rect 19432 24012 19484 24064
rect 20996 24157 21005 24191
rect 21005 24157 21039 24191
rect 21039 24157 21048 24191
rect 20996 24148 21048 24157
rect 21824 24148 21876 24200
rect 24676 24191 24728 24200
rect 20720 24080 20772 24132
rect 22100 24080 22152 24132
rect 23020 24012 23072 24064
rect 24676 24157 24685 24191
rect 24685 24157 24719 24191
rect 24719 24157 24728 24191
rect 24676 24148 24728 24157
rect 25228 24216 25280 24268
rect 27252 24216 27304 24268
rect 27988 24284 28040 24336
rect 30840 24352 30892 24404
rect 36728 24395 36780 24404
rect 36728 24361 36737 24395
rect 36737 24361 36771 24395
rect 36771 24361 36780 24395
rect 36728 24352 36780 24361
rect 25504 24148 25556 24200
rect 26792 24191 26844 24200
rect 26792 24157 26801 24191
rect 26801 24157 26835 24191
rect 26835 24157 26844 24191
rect 26792 24148 26844 24157
rect 27160 24148 27212 24200
rect 27528 24191 27580 24200
rect 27528 24157 27537 24191
rect 27537 24157 27571 24191
rect 27571 24157 27580 24191
rect 27528 24148 27580 24157
rect 28816 24148 28868 24200
rect 29644 24148 29696 24200
rect 26424 24080 26476 24132
rect 28540 24080 28592 24132
rect 32680 24284 32732 24336
rect 32496 24259 32548 24268
rect 32496 24225 32505 24259
rect 32505 24225 32539 24259
rect 32539 24225 32548 24259
rect 32496 24216 32548 24225
rect 33140 24216 33192 24268
rect 37280 24259 37332 24268
rect 30656 24148 30708 24200
rect 31024 24148 31076 24200
rect 32220 24191 32272 24200
rect 32220 24157 32229 24191
rect 32229 24157 32263 24191
rect 32263 24157 32272 24191
rect 32220 24148 32272 24157
rect 32312 24191 32364 24200
rect 32312 24157 32321 24191
rect 32321 24157 32355 24191
rect 32355 24157 32364 24191
rect 33232 24191 33284 24200
rect 32312 24148 32364 24157
rect 33232 24157 33241 24191
rect 33241 24157 33275 24191
rect 33275 24157 33284 24191
rect 33232 24148 33284 24157
rect 34704 24191 34756 24200
rect 34704 24157 34713 24191
rect 34713 24157 34747 24191
rect 34747 24157 34756 24191
rect 34704 24148 34756 24157
rect 34796 24148 34848 24200
rect 35348 24191 35400 24200
rect 35348 24157 35357 24191
rect 35357 24157 35391 24191
rect 35391 24157 35400 24191
rect 35348 24148 35400 24157
rect 37280 24225 37289 24259
rect 37289 24225 37323 24259
rect 37323 24225 37332 24259
rect 37280 24216 37332 24225
rect 37096 24148 37148 24200
rect 23480 24012 23532 24064
rect 24216 24012 24268 24064
rect 24308 24012 24360 24064
rect 25780 24012 25832 24064
rect 25964 24012 26016 24064
rect 28816 24055 28868 24064
rect 28816 24021 28825 24055
rect 28825 24021 28859 24055
rect 28859 24021 28868 24055
rect 28816 24012 28868 24021
rect 29644 24012 29696 24064
rect 31208 24012 31260 24064
rect 37280 24080 37332 24132
rect 32404 24012 32456 24064
rect 32956 24012 33008 24064
rect 34796 24055 34848 24064
rect 34796 24021 34805 24055
rect 34805 24021 34839 24055
rect 34839 24021 34848 24055
rect 34796 24012 34848 24021
rect 35624 24012 35676 24064
rect 37740 24055 37792 24064
rect 37740 24021 37749 24055
rect 37749 24021 37783 24055
rect 37783 24021 37792 24055
rect 37740 24012 37792 24021
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 11888 23851 11940 23860
rect 11888 23817 11897 23851
rect 11897 23817 11931 23851
rect 11931 23817 11940 23851
rect 11888 23808 11940 23817
rect 14280 23851 14332 23860
rect 14280 23817 14289 23851
rect 14289 23817 14323 23851
rect 14323 23817 14332 23851
rect 14280 23808 14332 23817
rect 15108 23808 15160 23860
rect 15936 23851 15988 23860
rect 15936 23817 15945 23851
rect 15945 23817 15979 23851
rect 15979 23817 15988 23851
rect 15936 23808 15988 23817
rect 17960 23851 18012 23860
rect 17960 23817 17969 23851
rect 17969 23817 18003 23851
rect 18003 23817 18012 23851
rect 17960 23808 18012 23817
rect 21364 23808 21416 23860
rect 22560 23808 22612 23860
rect 23848 23808 23900 23860
rect 24860 23808 24912 23860
rect 28080 23808 28132 23860
rect 29092 23851 29144 23860
rect 29092 23817 29101 23851
rect 29101 23817 29135 23851
rect 29135 23817 29144 23851
rect 29092 23808 29144 23817
rect 32312 23808 32364 23860
rect 33692 23808 33744 23860
rect 35348 23808 35400 23860
rect 35716 23808 35768 23860
rect 8576 23783 8628 23792
rect 8576 23749 8585 23783
rect 8585 23749 8619 23783
rect 8619 23749 8628 23783
rect 8576 23740 8628 23749
rect 10324 23740 10376 23792
rect 12716 23740 12768 23792
rect 14556 23740 14608 23792
rect 8392 23715 8444 23724
rect 8392 23681 8401 23715
rect 8401 23681 8435 23715
rect 8435 23681 8444 23715
rect 8392 23672 8444 23681
rect 9220 23715 9272 23724
rect 9220 23681 9229 23715
rect 9229 23681 9263 23715
rect 9263 23681 9272 23715
rect 9220 23672 9272 23681
rect 11152 23672 11204 23724
rect 12072 23715 12124 23724
rect 12072 23681 12081 23715
rect 12081 23681 12115 23715
rect 12115 23681 12124 23715
rect 12072 23672 12124 23681
rect 9312 23647 9364 23656
rect 9312 23613 9321 23647
rect 9321 23613 9355 23647
rect 9355 23613 9364 23647
rect 9312 23604 9364 23613
rect 10232 23604 10284 23656
rect 12532 23672 12584 23724
rect 10508 23536 10560 23588
rect 12348 23536 12400 23588
rect 13452 23715 13504 23724
rect 13452 23681 13461 23715
rect 13461 23681 13495 23715
rect 13495 23681 13504 23715
rect 13452 23672 13504 23681
rect 13636 23715 13688 23724
rect 13636 23681 13645 23715
rect 13645 23681 13679 23715
rect 13679 23681 13688 23715
rect 13636 23672 13688 23681
rect 14464 23715 14516 23724
rect 14464 23681 14473 23715
rect 14473 23681 14507 23715
rect 14507 23681 14516 23715
rect 14464 23672 14516 23681
rect 16396 23672 16448 23724
rect 18696 23740 18748 23792
rect 15200 23536 15252 23588
rect 16856 23604 16908 23656
rect 19432 23672 19484 23724
rect 21088 23715 21140 23724
rect 21088 23681 21097 23715
rect 21097 23681 21131 23715
rect 21131 23681 21140 23715
rect 21088 23672 21140 23681
rect 18604 23604 18656 23656
rect 18972 23647 19024 23656
rect 18972 23613 18981 23647
rect 18981 23613 19015 23647
rect 19015 23613 19024 23647
rect 18972 23604 19024 23613
rect 20444 23604 20496 23656
rect 22100 23715 22152 23724
rect 22100 23681 22109 23715
rect 22109 23681 22143 23715
rect 22143 23681 22152 23715
rect 22100 23672 22152 23681
rect 22744 23715 22796 23724
rect 22468 23604 22520 23656
rect 22744 23681 22753 23715
rect 22753 23681 22787 23715
rect 22787 23681 22796 23715
rect 22744 23672 22796 23681
rect 23480 23672 23532 23724
rect 23756 23672 23808 23724
rect 24952 23740 25004 23792
rect 29644 23783 29696 23792
rect 24400 23715 24452 23724
rect 24400 23681 24409 23715
rect 24409 23681 24443 23715
rect 24443 23681 24452 23715
rect 24400 23672 24452 23681
rect 25320 23604 25372 23656
rect 25688 23715 25740 23724
rect 25688 23681 25697 23715
rect 25697 23681 25731 23715
rect 25731 23681 25740 23715
rect 25688 23672 25740 23681
rect 26792 23672 26844 23724
rect 27252 23715 27304 23724
rect 27252 23681 27261 23715
rect 27261 23681 27295 23715
rect 27295 23681 27304 23715
rect 27252 23672 27304 23681
rect 27436 23715 27488 23724
rect 27436 23681 27445 23715
rect 27445 23681 27479 23715
rect 27479 23681 27488 23715
rect 27436 23672 27488 23681
rect 29644 23749 29653 23783
rect 29653 23749 29687 23783
rect 29687 23749 29696 23783
rect 29644 23740 29696 23749
rect 29828 23783 29880 23792
rect 29828 23749 29837 23783
rect 29837 23749 29871 23783
rect 29871 23749 29880 23783
rect 29828 23740 29880 23749
rect 32036 23740 32088 23792
rect 29276 23672 29328 23724
rect 30748 23672 30800 23724
rect 32680 23672 32732 23724
rect 33048 23715 33100 23724
rect 33048 23681 33057 23715
rect 33057 23681 33091 23715
rect 33091 23681 33100 23715
rect 33048 23672 33100 23681
rect 33600 23672 33652 23724
rect 35900 23740 35952 23792
rect 36636 23740 36688 23792
rect 29644 23604 29696 23656
rect 30656 23647 30708 23656
rect 30656 23613 30665 23647
rect 30665 23613 30699 23647
rect 30699 23613 30708 23647
rect 30656 23604 30708 23613
rect 33140 23604 33192 23656
rect 19984 23536 20036 23588
rect 23020 23536 23072 23588
rect 24952 23536 25004 23588
rect 26240 23536 26292 23588
rect 26976 23536 27028 23588
rect 27436 23536 27488 23588
rect 9680 23468 9732 23520
rect 10232 23511 10284 23520
rect 10232 23477 10241 23511
rect 10241 23477 10275 23511
rect 10275 23477 10284 23511
rect 10232 23468 10284 23477
rect 12808 23511 12860 23520
rect 12808 23477 12817 23511
rect 12817 23477 12851 23511
rect 12851 23477 12860 23511
rect 12808 23468 12860 23477
rect 13084 23468 13136 23520
rect 16488 23468 16540 23520
rect 17592 23468 17644 23520
rect 19340 23511 19392 23520
rect 19340 23477 19349 23511
rect 19349 23477 19383 23511
rect 19383 23477 19392 23511
rect 19340 23468 19392 23477
rect 26424 23468 26476 23520
rect 27160 23468 27212 23520
rect 27988 23511 28040 23520
rect 27988 23477 27997 23511
rect 27997 23477 28031 23511
rect 28031 23477 28040 23511
rect 27988 23468 28040 23477
rect 29000 23468 29052 23520
rect 33140 23511 33192 23520
rect 33140 23477 33149 23511
rect 33149 23477 33183 23511
rect 33183 23477 33192 23511
rect 33140 23468 33192 23477
rect 34612 23647 34664 23656
rect 34612 23613 34621 23647
rect 34621 23613 34655 23647
rect 34655 23613 34664 23647
rect 34612 23604 34664 23613
rect 35624 23604 35676 23656
rect 37188 23672 37240 23724
rect 37740 23604 37792 23656
rect 36728 23468 36780 23520
rect 37832 23511 37884 23520
rect 37832 23477 37841 23511
rect 37841 23477 37875 23511
rect 37875 23477 37884 23511
rect 37832 23468 37884 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 8392 23307 8444 23316
rect 8392 23273 8401 23307
rect 8401 23273 8435 23307
rect 8435 23273 8444 23307
rect 8392 23264 8444 23273
rect 9220 23264 9272 23316
rect 12532 23264 12584 23316
rect 15016 23264 15068 23316
rect 18788 23264 18840 23316
rect 10600 23196 10652 23248
rect 12256 23196 12308 23248
rect 9036 23128 9088 23180
rect 11152 23171 11204 23180
rect 11152 23137 11161 23171
rect 11161 23137 11195 23171
rect 11195 23137 11204 23171
rect 11152 23128 11204 23137
rect 11980 23128 12032 23180
rect 7012 23103 7064 23112
rect 7012 23069 7021 23103
rect 7021 23069 7055 23103
rect 7055 23069 7064 23103
rect 7012 23060 7064 23069
rect 8392 23060 8444 23112
rect 8944 23060 8996 23112
rect 10232 23103 10284 23112
rect 10232 23069 10241 23103
rect 10241 23069 10275 23103
rect 10275 23069 10284 23103
rect 10232 23060 10284 23069
rect 10416 23103 10468 23112
rect 10416 23069 10425 23103
rect 10425 23069 10459 23103
rect 10459 23069 10468 23103
rect 10416 23060 10468 23069
rect 10600 23103 10652 23112
rect 10600 23069 10609 23103
rect 10609 23069 10643 23103
rect 10643 23069 10652 23103
rect 10600 23060 10652 23069
rect 12716 23103 12768 23112
rect 11060 22924 11112 22976
rect 12716 23069 12725 23103
rect 12725 23069 12759 23103
rect 12759 23069 12768 23103
rect 12716 23060 12768 23069
rect 12900 23103 12952 23112
rect 12900 23069 12909 23103
rect 12909 23069 12943 23103
rect 12943 23069 12952 23103
rect 15108 23196 15160 23248
rect 17776 23239 17828 23248
rect 12900 23060 12952 23069
rect 13176 23060 13228 23112
rect 16764 23103 16816 23112
rect 16764 23069 16773 23103
rect 16773 23069 16807 23103
rect 16807 23069 16816 23103
rect 16764 23060 16816 23069
rect 17776 23205 17785 23239
rect 17785 23205 17819 23239
rect 17819 23205 17828 23239
rect 17776 23196 17828 23205
rect 17592 23103 17644 23112
rect 17592 23069 17601 23103
rect 17601 23069 17635 23103
rect 17635 23069 17644 23103
rect 17592 23060 17644 23069
rect 20260 23128 20312 23180
rect 20996 23264 21048 23316
rect 26608 23264 26660 23316
rect 26792 23307 26844 23316
rect 26792 23273 26801 23307
rect 26801 23273 26835 23307
rect 26835 23273 26844 23307
rect 26792 23264 26844 23273
rect 27804 23264 27856 23316
rect 28540 23307 28592 23316
rect 28540 23273 28549 23307
rect 28549 23273 28583 23307
rect 28583 23273 28592 23307
rect 28540 23264 28592 23273
rect 31484 23307 31536 23316
rect 21732 23196 21784 23248
rect 18788 23060 18840 23112
rect 19432 23103 19484 23112
rect 19432 23069 19441 23103
rect 19441 23069 19475 23103
rect 19475 23069 19484 23103
rect 19432 23060 19484 23069
rect 17960 22992 18012 23044
rect 20812 23060 20864 23112
rect 21548 23103 21600 23112
rect 21548 23069 21557 23103
rect 21557 23069 21591 23103
rect 21591 23069 21600 23103
rect 21548 23060 21600 23069
rect 24676 23196 24728 23248
rect 25688 23196 25740 23248
rect 23480 23060 23532 23112
rect 12624 22924 12676 22976
rect 14832 22924 14884 22976
rect 16396 22924 16448 22976
rect 22744 22992 22796 23044
rect 23756 23035 23808 23044
rect 23756 23001 23765 23035
rect 23765 23001 23799 23035
rect 23799 23001 23808 23035
rect 25044 23060 25096 23112
rect 25412 23103 25464 23112
rect 25412 23069 25421 23103
rect 25421 23069 25455 23103
rect 25455 23069 25464 23103
rect 25412 23060 25464 23069
rect 25872 23060 25924 23112
rect 26240 23060 26292 23112
rect 26608 23128 26660 23180
rect 27528 23128 27580 23180
rect 28080 23196 28132 23248
rect 28356 23128 28408 23180
rect 29000 23128 29052 23180
rect 23756 22992 23808 23001
rect 26884 23060 26936 23112
rect 27804 23103 27856 23112
rect 27068 22992 27120 23044
rect 27804 23069 27813 23103
rect 27813 23069 27847 23103
rect 27847 23069 27856 23103
rect 27804 23060 27856 23069
rect 27988 23060 28040 23112
rect 28816 23060 28868 23112
rect 29368 23128 29420 23180
rect 30380 23171 30432 23180
rect 30380 23137 30389 23171
rect 30389 23137 30423 23171
rect 30423 23137 30432 23171
rect 30380 23128 30432 23137
rect 31484 23273 31493 23307
rect 31493 23273 31527 23307
rect 31527 23273 31536 23307
rect 31484 23264 31536 23273
rect 33048 23264 33100 23316
rect 35624 23264 35676 23316
rect 36728 23307 36780 23316
rect 36728 23273 36737 23307
rect 36737 23273 36771 23307
rect 36771 23273 36780 23307
rect 36728 23264 36780 23273
rect 37096 23307 37148 23316
rect 37096 23273 37105 23307
rect 37105 23273 37139 23307
rect 37139 23273 37148 23307
rect 37096 23264 37148 23273
rect 37648 23307 37700 23316
rect 37648 23273 37657 23307
rect 37657 23273 37691 23307
rect 37691 23273 37700 23307
rect 37648 23264 37700 23273
rect 28632 22992 28684 23044
rect 32128 23196 32180 23248
rect 31944 23128 31996 23180
rect 31484 23103 31536 23112
rect 25688 22924 25740 22976
rect 26332 22924 26384 22976
rect 27252 22924 27304 22976
rect 31484 23069 31493 23103
rect 31493 23069 31527 23103
rect 31527 23069 31536 23103
rect 31484 23060 31536 23069
rect 33140 23060 33192 23112
rect 33692 23103 33744 23112
rect 33692 23069 33701 23103
rect 33701 23069 33735 23103
rect 33735 23069 33744 23103
rect 33692 23060 33744 23069
rect 35348 23060 35400 23112
rect 36636 23103 36688 23112
rect 36636 23069 36645 23103
rect 36645 23069 36679 23103
rect 36679 23069 36688 23103
rect 36636 23060 36688 23069
rect 37740 23060 37792 23112
rect 30840 22992 30892 23044
rect 32956 23035 33008 23044
rect 32956 23001 32965 23035
rect 32965 23001 32999 23035
rect 32999 23001 33008 23035
rect 32956 22992 33008 23001
rect 34796 22992 34848 23044
rect 35716 23035 35768 23044
rect 35716 23001 35725 23035
rect 35725 23001 35759 23035
rect 35759 23001 35768 23035
rect 35716 22992 35768 23001
rect 31024 22924 31076 22976
rect 33232 22924 33284 22976
rect 33416 22924 33468 22976
rect 33784 22967 33836 22976
rect 33784 22933 33793 22967
rect 33793 22933 33827 22967
rect 33827 22933 33836 22967
rect 33784 22924 33836 22933
rect 35440 22924 35492 22976
rect 35900 22967 35952 22976
rect 35900 22933 35925 22967
rect 35925 22933 35952 22967
rect 36084 22967 36136 22976
rect 35900 22924 35952 22933
rect 36084 22933 36093 22967
rect 36093 22933 36127 22967
rect 36127 22933 36136 22967
rect 36084 22924 36136 22933
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 9312 22720 9364 22772
rect 10416 22720 10468 22772
rect 12072 22720 12124 22772
rect 12900 22720 12952 22772
rect 16764 22720 16816 22772
rect 17684 22720 17736 22772
rect 14280 22695 14332 22704
rect 8944 22627 8996 22636
rect 8944 22593 8953 22627
rect 8953 22593 8987 22627
rect 8987 22593 8996 22627
rect 8944 22584 8996 22593
rect 9036 22627 9088 22636
rect 9036 22593 9045 22627
rect 9045 22593 9079 22627
rect 9079 22593 9088 22627
rect 9036 22584 9088 22593
rect 9864 22584 9916 22636
rect 10048 22627 10100 22636
rect 10048 22593 10057 22627
rect 10057 22593 10091 22627
rect 10091 22593 10100 22627
rect 10048 22584 10100 22593
rect 10508 22627 10560 22636
rect 10508 22593 10517 22627
rect 10517 22593 10551 22627
rect 10551 22593 10560 22627
rect 10508 22584 10560 22593
rect 11060 22584 11112 22636
rect 12072 22584 12124 22636
rect 12440 22584 12492 22636
rect 12808 22627 12860 22636
rect 12808 22593 12817 22627
rect 12817 22593 12851 22627
rect 12851 22593 12860 22627
rect 12808 22584 12860 22593
rect 14280 22661 14289 22695
rect 14289 22661 14323 22695
rect 14323 22661 14332 22695
rect 14280 22652 14332 22661
rect 14556 22652 14608 22704
rect 14832 22695 14884 22704
rect 14832 22661 14841 22695
rect 14841 22661 14875 22695
rect 14875 22661 14884 22695
rect 14832 22652 14884 22661
rect 8852 22559 8904 22568
rect 8852 22525 8861 22559
rect 8861 22525 8895 22559
rect 8895 22525 8904 22559
rect 8852 22516 8904 22525
rect 12348 22516 12400 22568
rect 12716 22516 12768 22568
rect 8760 22380 8812 22432
rect 9680 22380 9732 22432
rect 12072 22380 12124 22432
rect 13636 22516 13688 22568
rect 14372 22584 14424 22636
rect 15476 22584 15528 22636
rect 16396 22584 16448 22636
rect 18512 22652 18564 22704
rect 15660 22516 15712 22568
rect 15292 22448 15344 22500
rect 17040 22559 17092 22568
rect 17040 22525 17049 22559
rect 17049 22525 17083 22559
rect 17083 22525 17092 22559
rect 18604 22584 18656 22636
rect 19432 22720 19484 22772
rect 22652 22763 22704 22772
rect 22652 22729 22661 22763
rect 22661 22729 22695 22763
rect 22695 22729 22704 22763
rect 22652 22720 22704 22729
rect 23112 22720 23164 22772
rect 23204 22720 23256 22772
rect 23756 22720 23808 22772
rect 25044 22720 25096 22772
rect 24124 22652 24176 22704
rect 20260 22627 20312 22636
rect 20260 22593 20269 22627
rect 20269 22593 20303 22627
rect 20303 22593 20312 22627
rect 20260 22584 20312 22593
rect 20720 22584 20772 22636
rect 22744 22627 22796 22636
rect 22744 22593 22753 22627
rect 22753 22593 22787 22627
rect 22787 22593 22796 22627
rect 22744 22584 22796 22593
rect 23480 22627 23532 22636
rect 23480 22593 23489 22627
rect 23489 22593 23523 22627
rect 23523 22593 23532 22627
rect 23480 22584 23532 22593
rect 23572 22559 23624 22568
rect 17040 22516 17092 22525
rect 18052 22448 18104 22500
rect 22192 22448 22244 22500
rect 23572 22525 23581 22559
rect 23581 22525 23615 22559
rect 23615 22525 23624 22559
rect 23572 22516 23624 22525
rect 24584 22627 24636 22636
rect 24584 22593 24593 22627
rect 24593 22593 24627 22627
rect 24627 22593 24636 22627
rect 24768 22627 24820 22636
rect 24584 22584 24636 22593
rect 24768 22593 24777 22627
rect 24777 22593 24811 22627
rect 24811 22593 24820 22627
rect 24768 22584 24820 22593
rect 25228 22584 25280 22636
rect 25872 22720 25924 22772
rect 31024 22720 31076 22772
rect 27344 22695 27396 22704
rect 27344 22661 27353 22695
rect 27353 22661 27387 22695
rect 27387 22661 27396 22695
rect 27344 22652 27396 22661
rect 28724 22652 28776 22704
rect 26976 22627 27028 22636
rect 24308 22516 24360 22568
rect 26976 22593 26985 22627
rect 26985 22593 27019 22627
rect 27019 22593 27028 22627
rect 26976 22584 27028 22593
rect 27068 22627 27120 22636
rect 27068 22593 27078 22627
rect 27078 22593 27112 22627
rect 27112 22593 27120 22627
rect 27068 22584 27120 22593
rect 26884 22516 26936 22568
rect 27528 22584 27580 22636
rect 28540 22627 28592 22636
rect 27344 22516 27396 22568
rect 28540 22593 28549 22627
rect 28549 22593 28583 22627
rect 28583 22593 28592 22627
rect 28540 22584 28592 22593
rect 29092 22584 29144 22636
rect 29368 22627 29420 22636
rect 29000 22516 29052 22568
rect 29368 22593 29377 22627
rect 29377 22593 29411 22627
rect 29411 22593 29420 22627
rect 29368 22584 29420 22593
rect 30472 22584 30524 22636
rect 31944 22652 31996 22704
rect 30656 22516 30708 22568
rect 31392 22584 31444 22636
rect 33140 22720 33192 22772
rect 33600 22695 33652 22704
rect 32864 22584 32916 22636
rect 33600 22661 33609 22695
rect 33609 22661 33643 22695
rect 33643 22661 33652 22695
rect 33600 22652 33652 22661
rect 35624 22652 35676 22704
rect 36084 22627 36136 22636
rect 31484 22559 31536 22568
rect 31484 22525 31493 22559
rect 31493 22525 31527 22559
rect 31527 22525 31536 22559
rect 31484 22516 31536 22525
rect 33232 22516 33284 22568
rect 32128 22448 32180 22500
rect 15384 22380 15436 22432
rect 16488 22380 16540 22432
rect 20260 22380 20312 22432
rect 22008 22423 22060 22432
rect 22008 22389 22017 22423
rect 22017 22389 22051 22423
rect 22051 22389 22060 22423
rect 22008 22380 22060 22389
rect 22100 22380 22152 22432
rect 22652 22380 22704 22432
rect 25872 22380 25924 22432
rect 26792 22380 26844 22432
rect 27528 22380 27580 22432
rect 27804 22380 27856 22432
rect 28264 22380 28316 22432
rect 28724 22423 28776 22432
rect 28724 22389 28733 22423
rect 28733 22389 28767 22423
rect 28767 22389 28776 22423
rect 28724 22380 28776 22389
rect 29000 22380 29052 22432
rect 29920 22423 29972 22432
rect 29920 22389 29929 22423
rect 29929 22389 29963 22423
rect 29963 22389 29972 22423
rect 29920 22380 29972 22389
rect 33600 22448 33652 22500
rect 36084 22593 36093 22627
rect 36093 22593 36127 22627
rect 36127 22593 36136 22627
rect 36084 22584 36136 22593
rect 36268 22627 36320 22636
rect 36268 22593 36277 22627
rect 36277 22593 36311 22627
rect 36311 22593 36320 22627
rect 36268 22584 36320 22593
rect 33232 22380 33284 22432
rect 33968 22423 34020 22432
rect 33968 22389 33977 22423
rect 33977 22389 34011 22423
rect 34011 22389 34020 22423
rect 33968 22380 34020 22389
rect 34428 22423 34480 22432
rect 34428 22389 34437 22423
rect 34437 22389 34471 22423
rect 34471 22389 34480 22423
rect 34428 22380 34480 22389
rect 35532 22423 35584 22432
rect 35532 22389 35541 22423
rect 35541 22389 35575 22423
rect 35575 22389 35584 22423
rect 35900 22448 35952 22500
rect 36636 22448 36688 22500
rect 35532 22380 35584 22389
rect 36728 22380 36780 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 14464 22176 14516 22228
rect 11152 22151 11204 22160
rect 11152 22117 11161 22151
rect 11161 22117 11195 22151
rect 11195 22117 11204 22151
rect 11152 22108 11204 22117
rect 15200 22108 15252 22160
rect 15476 22151 15528 22160
rect 15476 22117 15485 22151
rect 15485 22117 15519 22151
rect 15519 22117 15528 22151
rect 15476 22108 15528 22117
rect 9680 22040 9732 22092
rect 9956 22083 10008 22092
rect 9956 22049 9965 22083
rect 9965 22049 9999 22083
rect 9999 22049 10008 22083
rect 9956 22040 10008 22049
rect 1400 22015 1452 22024
rect 1400 21981 1409 22015
rect 1409 21981 1443 22015
rect 1443 21981 1452 22015
rect 1400 21972 1452 21981
rect 8852 21972 8904 22024
rect 11612 21972 11664 22024
rect 10968 21947 11020 21956
rect 10968 21913 10977 21947
rect 10977 21913 11011 21947
rect 11011 21913 11020 21947
rect 10968 21904 11020 21913
rect 7932 21836 7984 21888
rect 11704 21836 11756 21888
rect 11977 22015 12029 22024
rect 11977 21981 12004 22015
rect 12004 21981 12029 22015
rect 11977 21972 12029 21981
rect 13084 22040 13136 22092
rect 17776 22176 17828 22228
rect 20720 22219 20772 22228
rect 20720 22185 20729 22219
rect 20729 22185 20763 22219
rect 20763 22185 20772 22219
rect 20720 22176 20772 22185
rect 22652 22219 22704 22228
rect 15660 22108 15712 22160
rect 22652 22185 22661 22219
rect 22661 22185 22695 22219
rect 22695 22185 22704 22219
rect 22652 22176 22704 22185
rect 22744 22176 22796 22228
rect 23664 22219 23716 22228
rect 23664 22185 23673 22219
rect 23673 22185 23707 22219
rect 23707 22185 23716 22219
rect 23664 22176 23716 22185
rect 25320 22176 25372 22228
rect 26056 22176 26108 22228
rect 26240 22219 26292 22228
rect 26240 22185 26249 22219
rect 26249 22185 26283 22219
rect 26283 22185 26292 22219
rect 26240 22176 26292 22185
rect 28172 22176 28224 22228
rect 28448 22176 28500 22228
rect 30564 22219 30616 22228
rect 16396 22083 16448 22092
rect 12256 22015 12308 22024
rect 12256 21981 12265 22015
rect 12265 21981 12299 22015
rect 12299 21981 12308 22015
rect 12256 21972 12308 21981
rect 14096 21972 14148 22024
rect 16396 22049 16405 22083
rect 16405 22049 16439 22083
rect 16439 22049 16448 22083
rect 16396 22040 16448 22049
rect 15200 21972 15252 22024
rect 15660 22015 15712 22024
rect 15384 21904 15436 21956
rect 15660 21981 15669 22015
rect 15669 21981 15703 22015
rect 15703 21981 15712 22015
rect 15660 21972 15712 21981
rect 15936 21972 15988 22024
rect 17776 22015 17828 22024
rect 17776 21981 17785 22015
rect 17785 21981 17819 22015
rect 17819 21981 17828 22015
rect 17776 21972 17828 21981
rect 18236 21972 18288 22024
rect 24400 22108 24452 22160
rect 24676 22108 24728 22160
rect 20352 22040 20404 22092
rect 23112 22083 23164 22092
rect 19064 21972 19116 22024
rect 19432 22015 19484 22024
rect 19432 21981 19441 22015
rect 19441 21981 19475 22015
rect 19475 21981 19484 22015
rect 19432 21972 19484 21981
rect 20260 22015 20312 22024
rect 20260 21981 20269 22015
rect 20269 21981 20303 22015
rect 20303 21981 20312 22015
rect 20260 21972 20312 21981
rect 23112 22049 23121 22083
rect 23121 22049 23155 22083
rect 23155 22049 23164 22083
rect 23112 22040 23164 22049
rect 16948 21904 17000 21956
rect 13084 21836 13136 21888
rect 13360 21879 13412 21888
rect 13360 21845 13369 21879
rect 13369 21845 13403 21879
rect 13403 21845 13412 21879
rect 13360 21836 13412 21845
rect 16304 21836 16356 21888
rect 17684 21947 17736 21956
rect 17684 21913 17693 21947
rect 17693 21913 17727 21947
rect 17727 21913 17736 21947
rect 17684 21904 17736 21913
rect 21548 21904 21600 21956
rect 22008 21904 22060 21956
rect 23664 22040 23716 22092
rect 23848 22083 23900 22092
rect 23848 22049 23857 22083
rect 23857 22049 23891 22083
rect 23891 22049 23900 22083
rect 24952 22083 25004 22092
rect 23848 22040 23900 22049
rect 23480 21972 23532 22024
rect 24952 22049 24961 22083
rect 24961 22049 24995 22083
rect 24995 22049 25004 22083
rect 24952 22040 25004 22049
rect 26516 22108 26568 22160
rect 26884 22108 26936 22160
rect 27712 22108 27764 22160
rect 28540 22108 28592 22160
rect 29828 22108 29880 22160
rect 30564 22185 30573 22219
rect 30573 22185 30607 22219
rect 30607 22185 30616 22219
rect 30564 22176 30616 22185
rect 34612 22176 34664 22228
rect 35624 22176 35676 22228
rect 33416 22108 33468 22160
rect 33692 22108 33744 22160
rect 33784 22108 33836 22160
rect 24584 21972 24636 22024
rect 24860 22015 24912 22024
rect 24860 21981 24869 22015
rect 24869 21981 24903 22015
rect 24903 21981 24912 22015
rect 24860 21972 24912 21981
rect 25412 21972 25464 22024
rect 27068 22040 27120 22092
rect 27528 22040 27580 22092
rect 28264 22083 28316 22092
rect 28264 22049 28273 22083
rect 28273 22049 28307 22083
rect 28307 22049 28316 22083
rect 28264 22040 28316 22049
rect 27988 21972 28040 22024
rect 29000 21972 29052 22024
rect 29552 22015 29604 22024
rect 29552 21981 29561 22015
rect 29561 21981 29595 22015
rect 29595 21981 29604 22015
rect 29552 21972 29604 21981
rect 29828 21972 29880 22024
rect 30748 22040 30800 22092
rect 31576 22040 31628 22092
rect 32496 22040 32548 22092
rect 31208 22015 31260 22024
rect 17132 21836 17184 21888
rect 18144 21836 18196 21888
rect 20812 21836 20864 21888
rect 21824 21879 21876 21888
rect 21824 21845 21833 21879
rect 21833 21845 21867 21879
rect 21867 21845 21876 21879
rect 21824 21836 21876 21845
rect 23480 21836 23532 21888
rect 26148 21836 26200 21888
rect 27160 21879 27212 21888
rect 27160 21845 27169 21879
rect 27169 21845 27203 21879
rect 27203 21845 27212 21879
rect 27160 21836 27212 21845
rect 27896 21879 27948 21888
rect 27896 21845 27905 21879
rect 27905 21845 27939 21879
rect 27939 21845 27948 21879
rect 27896 21836 27948 21845
rect 30656 21904 30708 21956
rect 28540 21836 28592 21888
rect 28724 21836 28776 21888
rect 30012 21836 30064 21888
rect 30104 21836 30156 21888
rect 31208 21981 31217 22015
rect 31217 21981 31251 22015
rect 31251 21981 31260 22015
rect 31208 21972 31260 21981
rect 32220 21972 32272 22024
rect 34060 21972 34112 22024
rect 35440 22015 35492 22024
rect 35440 21981 35449 22015
rect 35449 21981 35483 22015
rect 35483 21981 35492 22015
rect 35440 21972 35492 21981
rect 35624 22015 35676 22024
rect 35624 21981 35633 22015
rect 35633 21981 35667 22015
rect 35667 21981 35676 22015
rect 35624 21972 35676 21981
rect 37372 22015 37424 22024
rect 37372 21981 37381 22015
rect 37381 21981 37415 22015
rect 37415 21981 37424 22015
rect 37372 21972 37424 21981
rect 37740 22015 37792 22024
rect 37740 21981 37749 22015
rect 37749 21981 37783 22015
rect 37783 21981 37792 22015
rect 37740 21972 37792 21981
rect 30840 21836 30892 21888
rect 32496 21879 32548 21888
rect 32496 21845 32505 21879
rect 32505 21845 32539 21879
rect 32539 21845 32548 21879
rect 32496 21836 32548 21845
rect 34704 21879 34756 21888
rect 34704 21845 34713 21879
rect 34713 21845 34747 21879
rect 34747 21845 34756 21879
rect 34704 21836 34756 21845
rect 38108 21879 38160 21888
rect 38108 21845 38117 21879
rect 38117 21845 38151 21879
rect 38151 21845 38160 21879
rect 38108 21836 38160 21845
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 8852 21632 8904 21684
rect 10048 21632 10100 21684
rect 10232 21632 10284 21684
rect 9772 21564 9824 21616
rect 12624 21632 12676 21684
rect 13452 21632 13504 21684
rect 14372 21675 14424 21684
rect 14372 21641 14381 21675
rect 14381 21641 14415 21675
rect 14415 21641 14424 21675
rect 14372 21632 14424 21641
rect 7012 21428 7064 21480
rect 7288 21471 7340 21480
rect 7288 21437 7297 21471
rect 7297 21437 7331 21471
rect 7331 21437 7340 21471
rect 7288 21428 7340 21437
rect 11152 21428 11204 21480
rect 12624 21496 12676 21548
rect 13176 21564 13228 21616
rect 15384 21607 15436 21616
rect 15384 21573 15393 21607
rect 15393 21573 15427 21607
rect 15427 21573 15436 21607
rect 15384 21564 15436 21573
rect 13268 21539 13320 21548
rect 13268 21505 13302 21539
rect 13302 21505 13320 21539
rect 13268 21496 13320 21505
rect 15476 21496 15528 21548
rect 15936 21539 15988 21548
rect 15936 21505 15945 21539
rect 15945 21505 15979 21539
rect 15979 21505 15988 21539
rect 15936 21496 15988 21505
rect 16120 21539 16172 21548
rect 16120 21505 16129 21539
rect 16129 21505 16163 21539
rect 16163 21505 16172 21539
rect 16120 21496 16172 21505
rect 17316 21496 17368 21548
rect 20076 21675 20128 21684
rect 20076 21641 20085 21675
rect 20085 21641 20119 21675
rect 20119 21641 20128 21675
rect 20076 21632 20128 21641
rect 24032 21632 24084 21684
rect 22192 21564 22244 21616
rect 23388 21564 23440 21616
rect 23664 21564 23716 21616
rect 25412 21632 25464 21684
rect 18604 21539 18656 21548
rect 18604 21505 18613 21539
rect 18613 21505 18647 21539
rect 18647 21505 18656 21539
rect 18604 21496 18656 21505
rect 18880 21539 18932 21548
rect 18880 21505 18889 21539
rect 18889 21505 18923 21539
rect 18923 21505 18932 21539
rect 18880 21496 18932 21505
rect 19340 21496 19392 21548
rect 21824 21496 21876 21548
rect 22560 21539 22612 21548
rect 22560 21505 22569 21539
rect 22569 21505 22603 21539
rect 22603 21505 22612 21539
rect 22560 21496 22612 21505
rect 12808 21428 12860 21480
rect 14924 21428 14976 21480
rect 10140 21360 10192 21412
rect 12348 21403 12400 21412
rect 12348 21369 12357 21403
rect 12357 21369 12391 21403
rect 12391 21369 12400 21403
rect 12348 21360 12400 21369
rect 9864 21292 9916 21344
rect 12256 21292 12308 21344
rect 14372 21292 14424 21344
rect 15476 21292 15528 21344
rect 16580 21292 16632 21344
rect 23572 21496 23624 21548
rect 24400 21564 24452 21616
rect 24308 21539 24360 21548
rect 24308 21505 24317 21539
rect 24317 21505 24351 21539
rect 24351 21505 24360 21539
rect 24308 21496 24360 21505
rect 25228 21539 25280 21548
rect 23204 21360 23256 21412
rect 25228 21505 25237 21539
rect 25237 21505 25271 21539
rect 25271 21505 25280 21539
rect 25228 21496 25280 21505
rect 27896 21632 27948 21684
rect 27988 21632 28040 21684
rect 28540 21632 28592 21684
rect 28632 21632 28684 21684
rect 29000 21632 29052 21684
rect 29644 21675 29696 21684
rect 29644 21641 29653 21675
rect 29653 21641 29687 21675
rect 29687 21641 29696 21675
rect 29644 21632 29696 21641
rect 30012 21632 30064 21684
rect 32496 21632 32548 21684
rect 34060 21675 34112 21684
rect 34060 21641 34069 21675
rect 34069 21641 34103 21675
rect 34103 21641 34112 21675
rect 34060 21632 34112 21641
rect 37740 21632 37792 21684
rect 25872 21428 25924 21480
rect 26056 21539 26108 21548
rect 26056 21505 26065 21539
rect 26065 21505 26099 21539
rect 26099 21505 26108 21539
rect 26424 21564 26476 21616
rect 27068 21564 27120 21616
rect 29092 21564 29144 21616
rect 26056 21496 26108 21505
rect 26332 21539 26384 21548
rect 26332 21505 26341 21539
rect 26341 21505 26375 21539
rect 26375 21505 26384 21539
rect 26332 21496 26384 21505
rect 27344 21496 27396 21548
rect 28724 21539 28776 21548
rect 28724 21505 28733 21539
rect 28733 21505 28767 21539
rect 28767 21505 28776 21539
rect 28724 21496 28776 21505
rect 28908 21496 28960 21548
rect 29184 21496 29236 21548
rect 29368 21496 29420 21548
rect 29920 21564 29972 21616
rect 31576 21564 31628 21616
rect 30932 21496 30984 21548
rect 25228 21360 25280 21412
rect 26332 21360 26384 21412
rect 30564 21428 30616 21480
rect 20812 21335 20864 21344
rect 20812 21301 20821 21335
rect 20821 21301 20855 21335
rect 20855 21301 20864 21335
rect 20812 21292 20864 21301
rect 22284 21292 22336 21344
rect 23112 21292 23164 21344
rect 24124 21335 24176 21344
rect 24124 21301 24133 21335
rect 24133 21301 24167 21335
rect 24167 21301 24176 21335
rect 24124 21292 24176 21301
rect 24584 21292 24636 21344
rect 26056 21292 26108 21344
rect 26240 21292 26292 21344
rect 29552 21360 29604 21412
rect 30748 21360 30800 21412
rect 31300 21496 31352 21548
rect 32128 21539 32180 21548
rect 32128 21505 32137 21539
rect 32137 21505 32171 21539
rect 32171 21505 32180 21539
rect 32128 21496 32180 21505
rect 33968 21564 34020 21616
rect 34612 21564 34664 21616
rect 34704 21607 34756 21616
rect 34704 21573 34713 21607
rect 34713 21573 34747 21607
rect 34747 21573 34756 21607
rect 34704 21564 34756 21573
rect 34428 21496 34480 21548
rect 35532 21496 35584 21548
rect 35900 21539 35952 21548
rect 35900 21505 35909 21539
rect 35909 21505 35943 21539
rect 35943 21505 35952 21539
rect 35900 21496 35952 21505
rect 36084 21539 36136 21548
rect 36084 21505 36093 21539
rect 36093 21505 36127 21539
rect 36127 21505 36136 21539
rect 36084 21496 36136 21505
rect 35716 21428 35768 21480
rect 37648 21496 37700 21548
rect 37556 21471 37608 21480
rect 37556 21437 37565 21471
rect 37565 21437 37599 21471
rect 37599 21437 37608 21471
rect 37556 21428 37608 21437
rect 31208 21360 31260 21412
rect 35992 21360 36044 21412
rect 27896 21335 27948 21344
rect 27896 21301 27905 21335
rect 27905 21301 27939 21335
rect 27939 21301 27948 21335
rect 27896 21292 27948 21301
rect 28356 21292 28408 21344
rect 29644 21292 29696 21344
rect 30564 21292 30616 21344
rect 32404 21292 32456 21344
rect 34796 21292 34848 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 8576 21020 8628 21072
rect 9680 21088 9732 21140
rect 10140 21131 10192 21140
rect 10140 21097 10149 21131
rect 10149 21097 10183 21131
rect 10183 21097 10192 21131
rect 10140 21088 10192 21097
rect 9956 21020 10008 21072
rect 10416 21020 10468 21072
rect 10600 21020 10652 21072
rect 10048 20952 10100 21004
rect 10232 20952 10284 21004
rect 11796 21088 11848 21140
rect 12808 21131 12860 21140
rect 12808 21097 12817 21131
rect 12817 21097 12851 21131
rect 12851 21097 12860 21131
rect 12808 21088 12860 21097
rect 13084 21088 13136 21140
rect 16488 21088 16540 21140
rect 16948 21088 17000 21140
rect 13176 21020 13228 21072
rect 15660 21020 15712 21072
rect 16212 21020 16264 21072
rect 9772 20884 9824 20936
rect 10324 20884 10376 20936
rect 9864 20816 9916 20868
rect 10600 20927 10652 20936
rect 10600 20893 10609 20927
rect 10609 20893 10643 20927
rect 10643 20893 10652 20927
rect 13360 20952 13412 21004
rect 10600 20884 10652 20893
rect 11336 20884 11388 20936
rect 11704 20927 11756 20936
rect 11704 20893 11738 20927
rect 11738 20893 11756 20927
rect 11704 20884 11756 20893
rect 14372 20884 14424 20936
rect 17316 20952 17368 21004
rect 22560 21088 22612 21140
rect 27620 21088 27672 21140
rect 27712 21088 27764 21140
rect 33324 21131 33376 21140
rect 22192 21020 22244 21072
rect 23664 21020 23716 21072
rect 21640 20952 21692 21004
rect 11980 20816 12032 20868
rect 12808 20816 12860 20868
rect 13452 20816 13504 20868
rect 20076 20884 20128 20936
rect 21732 20884 21784 20936
rect 22468 20952 22520 21004
rect 23112 20884 23164 20936
rect 23477 20924 23529 20933
rect 23477 20890 23486 20924
rect 23486 20890 23520 20924
rect 23520 20890 23529 20924
rect 23477 20881 23529 20890
rect 23572 20927 23624 20936
rect 23572 20893 23581 20927
rect 23581 20893 23615 20927
rect 23615 20893 23624 20927
rect 24124 20952 24176 21004
rect 24952 20952 25004 21004
rect 25228 20952 25280 21004
rect 26332 20952 26384 21004
rect 27068 20952 27120 21004
rect 27896 20952 27948 21004
rect 28448 20952 28500 21004
rect 29644 20995 29696 21004
rect 23572 20884 23624 20893
rect 26792 20884 26844 20936
rect 28356 20927 28408 20936
rect 28356 20893 28365 20927
rect 28365 20893 28399 20927
rect 28399 20893 28408 20927
rect 28356 20884 28408 20893
rect 28540 20884 28592 20936
rect 28908 20884 28960 20936
rect 8392 20791 8444 20800
rect 8392 20757 8401 20791
rect 8401 20757 8435 20791
rect 8435 20757 8444 20791
rect 8392 20748 8444 20757
rect 9680 20791 9732 20800
rect 9680 20757 9689 20791
rect 9689 20757 9723 20791
rect 9723 20757 9732 20791
rect 9680 20748 9732 20757
rect 9772 20748 9824 20800
rect 10968 20748 11020 20800
rect 12624 20748 12676 20800
rect 13636 20748 13688 20800
rect 14280 20748 14332 20800
rect 15936 20748 15988 20800
rect 27896 20816 27948 20868
rect 20720 20748 20772 20800
rect 20904 20791 20956 20800
rect 20904 20757 20913 20791
rect 20913 20757 20947 20791
rect 20947 20757 20956 20791
rect 20904 20748 20956 20757
rect 23112 20791 23164 20800
rect 23112 20757 23121 20791
rect 23121 20757 23155 20791
rect 23155 20757 23164 20791
rect 23112 20748 23164 20757
rect 24860 20748 24912 20800
rect 25596 20748 25648 20800
rect 26424 20748 26476 20800
rect 28080 20859 28132 20868
rect 28080 20825 28089 20859
rect 28089 20825 28123 20859
rect 28123 20825 28132 20859
rect 28080 20816 28132 20825
rect 28448 20816 28500 20868
rect 29644 20961 29653 20995
rect 29653 20961 29687 20995
rect 29687 20961 29696 20995
rect 29644 20952 29696 20961
rect 33048 21020 33100 21072
rect 33324 21097 33333 21131
rect 33333 21097 33367 21131
rect 33367 21097 33376 21131
rect 33324 21088 33376 21097
rect 34888 21063 34940 21072
rect 34888 21029 34897 21063
rect 34897 21029 34931 21063
rect 34931 21029 34940 21063
rect 34888 21020 34940 21029
rect 31024 20995 31076 21004
rect 31024 20961 31033 20995
rect 31033 20961 31067 20995
rect 31067 20961 31076 20995
rect 31024 20952 31076 20961
rect 31576 20995 31628 21004
rect 31576 20961 31585 20995
rect 31585 20961 31619 20995
rect 31619 20961 31628 20995
rect 31576 20952 31628 20961
rect 34612 20952 34664 21004
rect 37648 21131 37700 21140
rect 37648 21097 37657 21131
rect 37657 21097 37691 21131
rect 37691 21097 37700 21131
rect 37648 21088 37700 21097
rect 35624 21020 35676 21072
rect 35900 21020 35952 21072
rect 35992 21020 36044 21072
rect 29276 20884 29328 20936
rect 30932 20927 30984 20936
rect 30932 20893 30941 20927
rect 30941 20893 30975 20927
rect 30975 20893 30984 20927
rect 30932 20884 30984 20893
rect 32128 20884 32180 20936
rect 32404 20927 32456 20936
rect 32404 20893 32413 20927
rect 32413 20893 32447 20927
rect 32447 20893 32456 20927
rect 32404 20884 32456 20893
rect 33232 20927 33284 20936
rect 33232 20893 33241 20927
rect 33241 20893 33275 20927
rect 33275 20893 33284 20927
rect 33232 20884 33284 20893
rect 34704 20927 34756 20936
rect 30748 20816 30800 20868
rect 32496 20816 32548 20868
rect 34704 20893 34713 20927
rect 34713 20893 34747 20927
rect 34747 20893 34756 20927
rect 34704 20884 34756 20893
rect 35532 20884 35584 20936
rect 35900 20927 35952 20936
rect 35900 20893 35909 20927
rect 35909 20893 35943 20927
rect 35943 20893 35952 20927
rect 35900 20884 35952 20893
rect 36084 20884 36136 20936
rect 37832 21020 37884 21072
rect 34888 20816 34940 20868
rect 29184 20748 29236 20800
rect 29368 20748 29420 20800
rect 31668 20748 31720 20800
rect 32036 20748 32088 20800
rect 33140 20748 33192 20800
rect 35440 20791 35492 20800
rect 35440 20757 35449 20791
rect 35449 20757 35483 20791
rect 35483 20757 35492 20791
rect 35440 20748 35492 20757
rect 35716 20748 35768 20800
rect 35900 20748 35952 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 10600 20544 10652 20596
rect 13268 20544 13320 20596
rect 14096 20544 14148 20596
rect 15292 20587 15344 20596
rect 15292 20553 15301 20587
rect 15301 20553 15335 20587
rect 15335 20553 15344 20587
rect 15292 20544 15344 20553
rect 17316 20587 17368 20596
rect 17316 20553 17325 20587
rect 17325 20553 17359 20587
rect 17359 20553 17368 20587
rect 17316 20544 17368 20553
rect 19432 20544 19484 20596
rect 20996 20544 21048 20596
rect 21732 20544 21784 20596
rect 21916 20544 21968 20596
rect 23572 20544 23624 20596
rect 8392 20408 8444 20460
rect 10048 20476 10100 20528
rect 7748 20340 7800 20392
rect 8760 20383 8812 20392
rect 8760 20349 8769 20383
rect 8769 20349 8803 20383
rect 8803 20349 8812 20383
rect 8760 20340 8812 20349
rect 9680 20408 9732 20460
rect 10324 20451 10376 20460
rect 10324 20417 10333 20451
rect 10333 20417 10367 20451
rect 10367 20417 10376 20451
rect 10324 20408 10376 20417
rect 10416 20451 10468 20460
rect 10416 20417 10425 20451
rect 10425 20417 10459 20451
rect 10459 20417 10468 20451
rect 10416 20408 10468 20417
rect 10968 20408 11020 20460
rect 12164 20383 12216 20392
rect 8300 20204 8352 20256
rect 12164 20349 12173 20383
rect 12173 20349 12207 20383
rect 12207 20349 12216 20383
rect 12164 20340 12216 20349
rect 13636 20383 13688 20392
rect 13636 20349 13645 20383
rect 13645 20349 13679 20383
rect 13679 20349 13688 20383
rect 13636 20340 13688 20349
rect 11980 20272 12032 20324
rect 14280 20451 14332 20460
rect 14280 20417 14289 20451
rect 14289 20417 14323 20451
rect 14323 20417 14332 20451
rect 14280 20408 14332 20417
rect 17868 20476 17920 20528
rect 18696 20476 18748 20528
rect 18972 20476 19024 20528
rect 20076 20476 20128 20528
rect 20720 20476 20772 20528
rect 17132 20408 17184 20460
rect 18052 20451 18104 20460
rect 18052 20417 18061 20451
rect 18061 20417 18095 20451
rect 18095 20417 18104 20451
rect 18052 20408 18104 20417
rect 15660 20340 15712 20392
rect 16396 20340 16448 20392
rect 17776 20340 17828 20392
rect 16580 20272 16632 20324
rect 20812 20408 20864 20460
rect 21180 20476 21232 20528
rect 22192 20476 22244 20528
rect 23664 20476 23716 20528
rect 24952 20519 25004 20528
rect 22008 20451 22060 20460
rect 22008 20417 22017 20451
rect 22017 20417 22051 20451
rect 22051 20417 22060 20451
rect 22008 20408 22060 20417
rect 22100 20451 22152 20460
rect 22100 20417 22109 20451
rect 22109 20417 22143 20451
rect 22143 20417 22152 20451
rect 22284 20451 22336 20460
rect 22100 20408 22152 20417
rect 22284 20417 22293 20451
rect 22293 20417 22327 20451
rect 22327 20417 22336 20451
rect 22284 20408 22336 20417
rect 22468 20451 22520 20460
rect 22468 20417 22477 20451
rect 22477 20417 22511 20451
rect 22511 20417 22520 20451
rect 22468 20408 22520 20417
rect 23020 20408 23072 20460
rect 23940 20451 23992 20460
rect 23940 20417 23949 20451
rect 23949 20417 23983 20451
rect 23983 20417 23992 20451
rect 23940 20408 23992 20417
rect 24216 20451 24268 20460
rect 24216 20417 24225 20451
rect 24225 20417 24259 20451
rect 24259 20417 24268 20451
rect 24216 20408 24268 20417
rect 24952 20485 24961 20519
rect 24961 20485 24995 20519
rect 24995 20485 25004 20519
rect 24952 20476 25004 20485
rect 25044 20408 25096 20460
rect 25780 20544 25832 20596
rect 29920 20544 29972 20596
rect 30932 20544 30984 20596
rect 26516 20476 26568 20528
rect 26792 20476 26844 20528
rect 26700 20408 26752 20460
rect 26884 20408 26936 20460
rect 27068 20451 27120 20460
rect 27068 20417 27077 20451
rect 27077 20417 27111 20451
rect 27111 20417 27120 20451
rect 27068 20408 27120 20417
rect 27712 20476 27764 20528
rect 27988 20476 28040 20528
rect 9128 20204 9180 20256
rect 15844 20204 15896 20256
rect 16856 20247 16908 20256
rect 16856 20213 16865 20247
rect 16865 20213 16899 20247
rect 16899 20213 16908 20247
rect 16856 20204 16908 20213
rect 20628 20272 20680 20324
rect 22836 20340 22888 20392
rect 23296 20340 23348 20392
rect 23480 20272 23532 20324
rect 25596 20272 25648 20324
rect 22376 20204 22428 20256
rect 25504 20204 25556 20256
rect 26332 20272 26384 20324
rect 28632 20408 28684 20460
rect 29000 20451 29052 20460
rect 29000 20417 29009 20451
rect 29009 20417 29043 20451
rect 29043 20417 29052 20451
rect 29000 20408 29052 20417
rect 29184 20476 29236 20528
rect 30104 20519 30156 20528
rect 30104 20485 30113 20519
rect 30113 20485 30147 20519
rect 30147 20485 30156 20519
rect 35440 20544 35492 20596
rect 30104 20476 30156 20485
rect 33232 20476 33284 20528
rect 28080 20340 28132 20392
rect 28724 20383 28776 20392
rect 28724 20349 28733 20383
rect 28733 20349 28767 20383
rect 28767 20349 28776 20383
rect 28724 20340 28776 20349
rect 32036 20408 32088 20460
rect 32128 20408 32180 20460
rect 32496 20451 32548 20460
rect 31668 20340 31720 20392
rect 32496 20417 32505 20451
rect 32505 20417 32539 20451
rect 32539 20417 32548 20451
rect 32496 20408 32548 20417
rect 33876 20476 33928 20528
rect 34796 20476 34848 20528
rect 33324 20340 33376 20392
rect 34704 20408 34756 20460
rect 36176 20451 36228 20460
rect 36176 20417 36185 20451
rect 36185 20417 36219 20451
rect 36219 20417 36228 20451
rect 36176 20408 36228 20417
rect 29184 20272 29236 20324
rect 35348 20340 35400 20392
rect 35992 20340 36044 20392
rect 26056 20247 26108 20256
rect 26056 20213 26065 20247
rect 26065 20213 26099 20247
rect 26099 20213 26108 20247
rect 26056 20204 26108 20213
rect 27712 20247 27764 20256
rect 27712 20213 27721 20247
rect 27721 20213 27755 20247
rect 27755 20213 27764 20247
rect 27712 20204 27764 20213
rect 31760 20204 31812 20256
rect 32588 20247 32640 20256
rect 32588 20213 32597 20247
rect 32597 20213 32631 20247
rect 32631 20213 32640 20247
rect 32588 20204 32640 20213
rect 32772 20204 32824 20256
rect 34244 20247 34296 20256
rect 34244 20213 34253 20247
rect 34253 20213 34287 20247
rect 34287 20213 34296 20247
rect 34244 20204 34296 20213
rect 35532 20204 35584 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 7748 20043 7800 20052
rect 7748 20009 7757 20043
rect 7757 20009 7791 20043
rect 7791 20009 7800 20043
rect 7748 20000 7800 20009
rect 7932 20000 7984 20052
rect 7932 19907 7984 19916
rect 7932 19873 7941 19907
rect 7941 19873 7975 19907
rect 7975 19873 7984 19907
rect 7932 19864 7984 19873
rect 9128 19932 9180 19984
rect 8392 19907 8444 19916
rect 8392 19873 8401 19907
rect 8401 19873 8435 19907
rect 8435 19873 8444 19907
rect 8392 19864 8444 19873
rect 10048 19932 10100 19984
rect 10968 19932 11020 19984
rect 8760 19796 8812 19848
rect 11980 19864 12032 19916
rect 12348 19907 12400 19916
rect 12348 19873 12357 19907
rect 12357 19873 12391 19907
rect 12391 19873 12400 19907
rect 12348 19864 12400 19873
rect 13452 19932 13504 19984
rect 12624 19907 12676 19916
rect 12624 19873 12633 19907
rect 12633 19873 12667 19907
rect 12667 19873 12676 19907
rect 12624 19864 12676 19873
rect 20076 20000 20128 20052
rect 22100 20000 22152 20052
rect 23664 20043 23716 20052
rect 23664 20009 23673 20043
rect 23673 20009 23707 20043
rect 23707 20009 23716 20043
rect 23664 20000 23716 20009
rect 24216 20000 24268 20052
rect 24768 20000 24820 20052
rect 17500 19932 17552 19984
rect 10416 19728 10468 19780
rect 11336 19796 11388 19848
rect 12808 19796 12860 19848
rect 14372 19839 14424 19848
rect 14372 19805 14381 19839
rect 14381 19805 14415 19839
rect 14415 19805 14424 19839
rect 14372 19796 14424 19805
rect 16120 19864 16172 19916
rect 16488 19907 16540 19916
rect 16488 19873 16497 19907
rect 16497 19873 16531 19907
rect 16531 19873 16540 19907
rect 16488 19864 16540 19873
rect 17868 19907 17920 19916
rect 17868 19873 17877 19907
rect 17877 19873 17911 19907
rect 17911 19873 17920 19907
rect 17868 19864 17920 19873
rect 18236 19864 18288 19916
rect 15844 19796 15896 19848
rect 17960 19796 18012 19848
rect 19984 19839 20036 19848
rect 10508 19703 10560 19712
rect 10508 19669 10517 19703
rect 10517 19669 10551 19703
rect 10551 19669 10560 19703
rect 10508 19660 10560 19669
rect 10600 19660 10652 19712
rect 14280 19728 14332 19780
rect 19340 19771 19392 19780
rect 19340 19737 19349 19771
rect 19349 19737 19383 19771
rect 19383 19737 19392 19771
rect 19340 19728 19392 19737
rect 19984 19805 19993 19839
rect 19993 19805 20027 19839
rect 20027 19805 20036 19839
rect 19984 19796 20036 19805
rect 20628 19796 20680 19848
rect 26148 19932 26200 19984
rect 26884 19975 26936 19984
rect 20996 19907 21048 19916
rect 20996 19873 21005 19907
rect 21005 19873 21039 19907
rect 21039 19873 21048 19907
rect 20996 19864 21048 19873
rect 22192 19864 22244 19916
rect 23848 19907 23900 19916
rect 21180 19796 21232 19848
rect 22376 19796 22428 19848
rect 23848 19873 23857 19907
rect 23857 19873 23891 19907
rect 23891 19873 23900 19907
rect 23848 19864 23900 19873
rect 24768 19907 24820 19916
rect 24768 19873 24777 19907
rect 24777 19873 24811 19907
rect 24811 19873 24820 19907
rect 24768 19864 24820 19873
rect 25780 19864 25832 19916
rect 26884 19941 26893 19975
rect 26893 19941 26927 19975
rect 26927 19941 26936 19975
rect 26884 19932 26936 19941
rect 28356 20000 28408 20052
rect 28724 20000 28776 20052
rect 32128 20000 32180 20052
rect 32772 20043 32824 20052
rect 32772 20009 32781 20043
rect 32781 20009 32815 20043
rect 32815 20009 32824 20043
rect 32772 20000 32824 20009
rect 36176 20000 36228 20052
rect 29276 19932 29328 19984
rect 22836 19839 22888 19848
rect 22836 19805 22845 19839
rect 22845 19805 22879 19839
rect 22879 19805 22888 19839
rect 22836 19796 22888 19805
rect 23388 19796 23440 19848
rect 23572 19839 23624 19848
rect 23572 19805 23581 19839
rect 23581 19805 23615 19839
rect 23615 19805 23624 19839
rect 23572 19796 23624 19805
rect 23940 19796 23992 19848
rect 24492 19796 24544 19848
rect 20168 19771 20220 19780
rect 20168 19737 20177 19771
rect 20177 19737 20211 19771
rect 20211 19737 20220 19771
rect 20168 19728 20220 19737
rect 22652 19771 22704 19780
rect 11060 19660 11112 19712
rect 12624 19660 12676 19712
rect 13452 19703 13504 19712
rect 13452 19669 13461 19703
rect 13461 19669 13495 19703
rect 13495 19669 13504 19703
rect 13452 19660 13504 19669
rect 15660 19660 15712 19712
rect 20536 19660 20588 19712
rect 22652 19737 22661 19771
rect 22661 19737 22695 19771
rect 22695 19737 22704 19771
rect 22652 19728 22704 19737
rect 22744 19771 22796 19780
rect 22744 19737 22753 19771
rect 22753 19737 22787 19771
rect 22787 19737 22796 19771
rect 22744 19728 22796 19737
rect 22928 19728 22980 19780
rect 24860 19839 24912 19848
rect 24860 19805 24869 19839
rect 24869 19805 24903 19839
rect 24903 19805 24912 19839
rect 24860 19796 24912 19805
rect 25044 19839 25096 19848
rect 25044 19805 25053 19839
rect 25053 19805 25087 19839
rect 25087 19805 25096 19839
rect 25044 19796 25096 19805
rect 25964 19796 26016 19848
rect 26332 19796 26384 19848
rect 28448 19796 28500 19848
rect 29000 19796 29052 19848
rect 29368 19796 29420 19848
rect 29736 19839 29788 19848
rect 29736 19805 29745 19839
rect 29745 19805 29779 19839
rect 29779 19805 29788 19839
rect 29736 19796 29788 19805
rect 30564 19839 30616 19848
rect 30564 19805 30573 19839
rect 30573 19805 30607 19839
rect 30607 19805 30616 19839
rect 30564 19796 30616 19805
rect 31116 19796 31168 19848
rect 32036 19864 32088 19916
rect 31668 19839 31720 19848
rect 31668 19805 31677 19839
rect 31677 19805 31711 19839
rect 31711 19805 31720 19839
rect 31668 19796 31720 19805
rect 34796 19932 34848 19984
rect 34244 19864 34296 19916
rect 35256 19864 35308 19916
rect 35348 19796 35400 19848
rect 28908 19728 28960 19780
rect 34336 19728 34388 19780
rect 23020 19703 23072 19712
rect 23020 19669 23029 19703
rect 23029 19669 23063 19703
rect 23063 19669 23072 19703
rect 23020 19660 23072 19669
rect 23480 19660 23532 19712
rect 25780 19660 25832 19712
rect 26516 19660 26568 19712
rect 28172 19660 28224 19712
rect 28448 19703 28500 19712
rect 28448 19669 28457 19703
rect 28457 19669 28491 19703
rect 28491 19669 28500 19703
rect 28448 19660 28500 19669
rect 29552 19660 29604 19712
rect 30472 19660 30524 19712
rect 31024 19660 31076 19712
rect 32404 19703 32456 19712
rect 32404 19669 32413 19703
rect 32413 19669 32447 19703
rect 32447 19669 32456 19703
rect 32404 19660 32456 19669
rect 33048 19660 33100 19712
rect 34980 19660 35032 19712
rect 35440 19660 35492 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 9128 19499 9180 19508
rect 9128 19465 9137 19499
rect 9137 19465 9171 19499
rect 9171 19465 9180 19499
rect 9128 19456 9180 19465
rect 10324 19456 10376 19508
rect 7288 19388 7340 19440
rect 9404 19388 9456 19440
rect 10232 19388 10284 19440
rect 15936 19456 15988 19508
rect 16488 19456 16540 19508
rect 17132 19456 17184 19508
rect 19984 19456 20036 19508
rect 8024 19363 8076 19372
rect 8024 19329 8058 19363
rect 8058 19329 8076 19363
rect 10324 19363 10376 19372
rect 8024 19320 8076 19329
rect 10324 19329 10333 19363
rect 10333 19329 10367 19363
rect 10367 19329 10376 19363
rect 10324 19320 10376 19329
rect 10600 19388 10652 19440
rect 10784 19388 10836 19440
rect 10968 19388 11020 19440
rect 11980 19388 12032 19440
rect 12348 19388 12400 19440
rect 19800 19388 19852 19440
rect 13452 19363 13504 19372
rect 13452 19329 13461 19363
rect 13461 19329 13495 19363
rect 13495 19329 13504 19363
rect 13452 19320 13504 19329
rect 13636 19363 13688 19372
rect 13636 19329 13645 19363
rect 13645 19329 13679 19363
rect 13679 19329 13688 19363
rect 13636 19320 13688 19329
rect 10600 19295 10652 19304
rect 10600 19261 10609 19295
rect 10609 19261 10643 19295
rect 10643 19261 10652 19295
rect 10600 19252 10652 19261
rect 12256 19295 12308 19304
rect 12256 19261 12265 19295
rect 12265 19261 12299 19295
rect 12299 19261 12308 19295
rect 12256 19252 12308 19261
rect 12716 19252 12768 19304
rect 10784 19184 10836 19236
rect 12440 19184 12492 19236
rect 13176 19252 13228 19304
rect 13820 19320 13872 19372
rect 15384 19363 15436 19372
rect 15384 19329 15393 19363
rect 15393 19329 15427 19363
rect 15427 19329 15436 19363
rect 15384 19320 15436 19329
rect 16948 19363 17000 19372
rect 16948 19329 16957 19363
rect 16957 19329 16991 19363
rect 16991 19329 17000 19363
rect 16948 19320 17000 19329
rect 17224 19363 17276 19372
rect 17224 19329 17258 19363
rect 17258 19329 17276 19363
rect 17224 19320 17276 19329
rect 18788 19320 18840 19372
rect 15660 19295 15712 19304
rect 15660 19261 15669 19295
rect 15669 19261 15703 19295
rect 15703 19261 15712 19295
rect 15660 19252 15712 19261
rect 19248 19363 19300 19372
rect 19248 19329 19257 19363
rect 19257 19329 19291 19363
rect 19291 19329 19300 19363
rect 20352 19456 20404 19508
rect 21088 19456 21140 19508
rect 22744 19456 22796 19508
rect 25596 19499 25648 19508
rect 25596 19465 25605 19499
rect 25605 19465 25639 19499
rect 25639 19465 25648 19499
rect 25596 19456 25648 19465
rect 20904 19388 20956 19440
rect 19248 19320 19300 19329
rect 19156 19252 19208 19304
rect 19800 19252 19852 19304
rect 12624 19159 12676 19168
rect 12624 19125 12633 19159
rect 12633 19125 12667 19159
rect 12667 19125 12676 19159
rect 12624 19116 12676 19125
rect 12992 19116 13044 19168
rect 13360 19116 13412 19168
rect 16764 19184 16816 19236
rect 15016 19159 15068 19168
rect 15016 19125 15025 19159
rect 15025 19125 15059 19159
rect 15059 19125 15068 19159
rect 15016 19116 15068 19125
rect 15108 19116 15160 19168
rect 20536 19320 20588 19372
rect 22652 19388 22704 19440
rect 20352 19252 20404 19304
rect 23756 19320 23808 19372
rect 23848 19320 23900 19372
rect 25504 19320 25556 19372
rect 25596 19320 25648 19372
rect 26240 19456 26292 19508
rect 27344 19388 27396 19440
rect 29644 19431 29696 19440
rect 29644 19397 29653 19431
rect 29653 19397 29687 19431
rect 29687 19397 29696 19431
rect 29644 19388 29696 19397
rect 29920 19456 29972 19508
rect 33876 19499 33928 19508
rect 33876 19465 33885 19499
rect 33885 19465 33919 19499
rect 33919 19465 33928 19499
rect 33876 19456 33928 19465
rect 34980 19456 35032 19508
rect 30564 19388 30616 19440
rect 31116 19388 31168 19440
rect 32588 19388 32640 19440
rect 32864 19388 32916 19440
rect 25780 19363 25832 19372
rect 25780 19329 25789 19363
rect 25789 19329 25823 19363
rect 25823 19329 25832 19363
rect 25780 19320 25832 19329
rect 26240 19363 26292 19372
rect 21916 19252 21968 19304
rect 24492 19252 24544 19304
rect 26240 19329 26249 19363
rect 26249 19329 26283 19363
rect 26283 19329 26292 19363
rect 26240 19320 26292 19329
rect 28448 19320 28500 19372
rect 29000 19320 29052 19372
rect 29552 19363 29604 19372
rect 29552 19329 29561 19363
rect 29561 19329 29595 19363
rect 29595 19329 29604 19363
rect 29552 19320 29604 19329
rect 20536 19184 20588 19236
rect 20996 19184 21048 19236
rect 23572 19184 23624 19236
rect 25780 19184 25832 19236
rect 26056 19252 26108 19304
rect 32128 19363 32180 19372
rect 32128 19329 32137 19363
rect 32137 19329 32171 19363
rect 32171 19329 32180 19363
rect 32128 19320 32180 19329
rect 27896 19184 27948 19236
rect 20260 19116 20312 19168
rect 20812 19116 20864 19168
rect 23296 19116 23348 19168
rect 25688 19116 25740 19168
rect 26056 19116 26108 19168
rect 26240 19116 26292 19168
rect 30196 19252 30248 19304
rect 31760 19252 31812 19304
rect 32680 19320 32732 19372
rect 35348 19388 35400 19440
rect 34060 19363 34112 19372
rect 34060 19329 34069 19363
rect 34069 19329 34103 19363
rect 34103 19329 34112 19363
rect 34060 19320 34112 19329
rect 34152 19363 34204 19372
rect 34152 19329 34161 19363
rect 34161 19329 34195 19363
rect 34195 19329 34204 19363
rect 34152 19320 34204 19329
rect 34612 19320 34664 19372
rect 28724 19184 28776 19236
rect 32404 19184 32456 19236
rect 33140 19184 33192 19236
rect 34704 19252 34756 19304
rect 34796 19184 34848 19236
rect 29092 19116 29144 19168
rect 29368 19159 29420 19168
rect 29368 19125 29377 19159
rect 29377 19125 29411 19159
rect 29411 19125 29420 19159
rect 29368 19116 29420 19125
rect 31116 19116 31168 19168
rect 31300 19116 31352 19168
rect 33968 19116 34020 19168
rect 35532 19116 35584 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 8024 18912 8076 18964
rect 10324 18912 10376 18964
rect 10600 18912 10652 18964
rect 13820 18912 13872 18964
rect 13912 18912 13964 18964
rect 15108 18912 15160 18964
rect 15384 18912 15436 18964
rect 16764 18912 16816 18964
rect 10232 18819 10284 18828
rect 10232 18785 10241 18819
rect 10241 18785 10275 18819
rect 10275 18785 10284 18819
rect 10232 18776 10284 18785
rect 8300 18751 8352 18760
rect 8300 18717 8309 18751
rect 8309 18717 8343 18751
rect 8343 18717 8352 18751
rect 8300 18708 8352 18717
rect 9680 18751 9732 18760
rect 9680 18717 9689 18751
rect 9689 18717 9723 18751
rect 9723 18717 9732 18751
rect 9680 18708 9732 18717
rect 10416 18708 10468 18760
rect 11888 18708 11940 18760
rect 14372 18751 14424 18760
rect 14372 18717 14381 18751
rect 14381 18717 14415 18751
rect 14415 18717 14424 18751
rect 16948 18776 17000 18828
rect 16396 18751 16448 18760
rect 14372 18708 14424 18717
rect 16396 18717 16405 18751
rect 16405 18717 16439 18751
rect 16439 18717 16448 18751
rect 16396 18708 16448 18717
rect 19340 18912 19392 18964
rect 22008 18912 22060 18964
rect 23572 18912 23624 18964
rect 23848 18955 23900 18964
rect 23848 18921 23857 18955
rect 23857 18921 23891 18955
rect 23891 18921 23900 18955
rect 23848 18912 23900 18921
rect 24860 18912 24912 18964
rect 27896 18912 27948 18964
rect 29276 18912 29328 18964
rect 17960 18844 18012 18896
rect 18696 18844 18748 18896
rect 23296 18844 23348 18896
rect 18420 18776 18472 18828
rect 20904 18776 20956 18828
rect 24676 18844 24728 18896
rect 29368 18844 29420 18896
rect 24308 18776 24360 18828
rect 30472 18912 30524 18964
rect 31760 18955 31812 18964
rect 31760 18921 31769 18955
rect 31769 18921 31803 18955
rect 31803 18921 31812 18955
rect 31760 18912 31812 18921
rect 34060 18844 34112 18896
rect 34520 18776 34572 18828
rect 34980 18819 35032 18828
rect 34980 18785 34989 18819
rect 34989 18785 35023 18819
rect 35023 18785 35032 18819
rect 34980 18776 35032 18785
rect 18236 18751 18288 18760
rect 18236 18717 18245 18751
rect 18245 18717 18279 18751
rect 18279 18717 18288 18751
rect 18236 18708 18288 18717
rect 19708 18751 19760 18760
rect 19708 18717 19717 18751
rect 19717 18717 19751 18751
rect 19751 18717 19760 18751
rect 19708 18708 19760 18717
rect 21916 18751 21968 18760
rect 21916 18717 21925 18751
rect 21925 18717 21959 18751
rect 21959 18717 21968 18751
rect 21916 18708 21968 18717
rect 23112 18708 23164 18760
rect 24492 18708 24544 18760
rect 25044 18751 25096 18760
rect 9772 18640 9824 18692
rect 12716 18640 12768 18692
rect 16304 18640 16356 18692
rect 16580 18683 16632 18692
rect 16580 18649 16589 18683
rect 16589 18649 16623 18683
rect 16623 18649 16632 18683
rect 16580 18640 16632 18649
rect 16764 18640 16816 18692
rect 18144 18683 18196 18692
rect 18144 18649 18153 18683
rect 18153 18649 18187 18683
rect 18187 18649 18196 18683
rect 18144 18640 18196 18649
rect 24124 18640 24176 18692
rect 11244 18572 11296 18624
rect 17960 18572 18012 18624
rect 18972 18572 19024 18624
rect 21824 18572 21876 18624
rect 21916 18572 21968 18624
rect 22744 18572 22796 18624
rect 23296 18572 23348 18624
rect 23572 18572 23624 18624
rect 25044 18717 25053 18751
rect 25053 18717 25087 18751
rect 25087 18717 25096 18751
rect 25044 18708 25096 18717
rect 25504 18751 25556 18760
rect 25504 18717 25513 18751
rect 25513 18717 25547 18751
rect 25547 18717 25556 18751
rect 25504 18708 25556 18717
rect 25872 18751 25924 18760
rect 25872 18717 25881 18751
rect 25881 18717 25915 18751
rect 25915 18717 25924 18751
rect 25872 18708 25924 18717
rect 26332 18708 26384 18760
rect 26792 18751 26844 18760
rect 26792 18717 26801 18751
rect 26801 18717 26835 18751
rect 26835 18717 26844 18751
rect 26792 18708 26844 18717
rect 26976 18708 27028 18760
rect 26240 18640 26292 18692
rect 29460 18708 29512 18760
rect 29736 18751 29788 18760
rect 29736 18717 29745 18751
rect 29745 18717 29779 18751
rect 29779 18717 29788 18751
rect 29736 18708 29788 18717
rect 29920 18751 29972 18760
rect 29920 18717 29929 18751
rect 29929 18717 29963 18751
rect 29963 18717 29972 18751
rect 29920 18708 29972 18717
rect 30196 18751 30248 18760
rect 30196 18717 30205 18751
rect 30205 18717 30239 18751
rect 30239 18717 30248 18751
rect 30196 18708 30248 18717
rect 30840 18751 30892 18760
rect 30840 18717 30849 18751
rect 30849 18717 30883 18751
rect 30883 18717 30892 18751
rect 30840 18708 30892 18717
rect 31024 18708 31076 18760
rect 31668 18708 31720 18760
rect 31852 18751 31904 18760
rect 31852 18717 31861 18751
rect 31861 18717 31895 18751
rect 31895 18717 31904 18751
rect 32680 18751 32732 18760
rect 31852 18708 31904 18717
rect 32680 18717 32689 18751
rect 32689 18717 32723 18751
rect 32723 18717 32732 18751
rect 32680 18708 32732 18717
rect 32864 18708 32916 18760
rect 33140 18751 33192 18760
rect 33140 18717 33149 18751
rect 33149 18717 33183 18751
rect 33183 18717 33192 18751
rect 33140 18708 33192 18717
rect 33968 18751 34020 18760
rect 33968 18717 33977 18751
rect 33977 18717 34011 18751
rect 34011 18717 34020 18751
rect 33968 18708 34020 18717
rect 34796 18708 34848 18760
rect 25136 18572 25188 18624
rect 26148 18572 26200 18624
rect 26976 18615 27028 18624
rect 26976 18581 26985 18615
rect 26985 18581 27019 18615
rect 27019 18581 27028 18615
rect 26976 18572 27028 18581
rect 28724 18572 28776 18624
rect 30104 18640 30156 18692
rect 33232 18640 33284 18692
rect 31116 18572 31168 18624
rect 32404 18572 32456 18624
rect 32956 18572 33008 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 12716 18411 12768 18420
rect 12716 18377 12725 18411
rect 12725 18377 12759 18411
rect 12759 18377 12768 18411
rect 12716 18368 12768 18377
rect 14004 18411 14056 18420
rect 10508 18300 10560 18352
rect 9404 18275 9456 18284
rect 9404 18241 9413 18275
rect 9413 18241 9447 18275
rect 9447 18241 9456 18275
rect 9404 18232 9456 18241
rect 11888 18232 11940 18284
rect 10784 18139 10836 18148
rect 10784 18105 10793 18139
rect 10793 18105 10827 18139
rect 10827 18105 10836 18139
rect 12440 18300 12492 18352
rect 12992 18232 13044 18284
rect 13176 18275 13228 18284
rect 13176 18241 13185 18275
rect 13185 18241 13219 18275
rect 13219 18241 13228 18275
rect 13176 18232 13228 18241
rect 14004 18377 14013 18411
rect 14013 18377 14047 18411
rect 14047 18377 14056 18411
rect 14004 18368 14056 18377
rect 16580 18368 16632 18420
rect 16948 18368 17000 18420
rect 18144 18368 18196 18420
rect 23664 18368 23716 18420
rect 25596 18411 25648 18420
rect 25596 18377 25605 18411
rect 25605 18377 25639 18411
rect 25639 18377 25648 18411
rect 25596 18368 25648 18377
rect 25872 18368 25924 18420
rect 26976 18368 27028 18420
rect 29736 18368 29788 18420
rect 31208 18368 31260 18420
rect 32680 18368 32732 18420
rect 33232 18368 33284 18420
rect 13820 18300 13872 18352
rect 15936 18343 15988 18352
rect 15936 18309 15945 18343
rect 15945 18309 15979 18343
rect 15979 18309 15988 18343
rect 15936 18300 15988 18309
rect 17040 18343 17092 18352
rect 17040 18309 17049 18343
rect 17049 18309 17083 18343
rect 17083 18309 17092 18343
rect 17040 18300 17092 18309
rect 17132 18343 17184 18352
rect 17132 18309 17141 18343
rect 17141 18309 17175 18343
rect 17175 18309 17184 18343
rect 17132 18300 17184 18309
rect 19340 18300 19392 18352
rect 15292 18275 15344 18284
rect 10784 18096 10836 18105
rect 15292 18241 15301 18275
rect 15301 18241 15335 18275
rect 15335 18241 15344 18275
rect 15292 18232 15344 18241
rect 16488 18232 16540 18284
rect 16396 18164 16448 18216
rect 17040 18164 17092 18216
rect 18236 18232 18288 18284
rect 19248 18232 19300 18284
rect 20168 18232 20220 18284
rect 23480 18300 23532 18352
rect 21824 18275 21876 18284
rect 21824 18241 21833 18275
rect 21833 18241 21867 18275
rect 21867 18241 21876 18275
rect 21824 18232 21876 18241
rect 22008 18275 22060 18284
rect 22008 18241 22017 18275
rect 22017 18241 22051 18275
rect 22051 18241 22060 18275
rect 22008 18232 22060 18241
rect 23572 18232 23624 18284
rect 24768 18232 24820 18284
rect 25964 18300 26016 18352
rect 26792 18300 26844 18352
rect 25780 18232 25832 18284
rect 26148 18275 26200 18284
rect 26148 18241 26157 18275
rect 26157 18241 26191 18275
rect 26191 18241 26200 18275
rect 26148 18232 26200 18241
rect 22744 18207 22796 18216
rect 22744 18173 22753 18207
rect 22753 18173 22787 18207
rect 22787 18173 22796 18207
rect 22744 18164 22796 18173
rect 25320 18164 25372 18216
rect 16764 18096 16816 18148
rect 17224 18096 17276 18148
rect 26056 18096 26108 18148
rect 30196 18300 30248 18352
rect 28724 18275 28776 18284
rect 28724 18241 28733 18275
rect 28733 18241 28767 18275
rect 28767 18241 28776 18275
rect 28724 18232 28776 18241
rect 31392 18300 31444 18352
rect 32404 18300 32456 18352
rect 31300 18232 31352 18284
rect 31668 18232 31720 18284
rect 32128 18275 32180 18284
rect 32128 18241 32137 18275
rect 32137 18241 32171 18275
rect 32171 18241 32180 18275
rect 32128 18232 32180 18241
rect 32956 18275 33008 18284
rect 32956 18241 32965 18275
rect 32965 18241 32999 18275
rect 32999 18241 33008 18275
rect 32956 18232 33008 18241
rect 33968 18368 34020 18420
rect 34980 18411 35032 18420
rect 34980 18377 34989 18411
rect 34989 18377 35023 18411
rect 35023 18377 35032 18411
rect 34980 18368 35032 18377
rect 34152 18232 34204 18284
rect 35348 18232 35400 18284
rect 31116 18164 31168 18216
rect 31484 18164 31536 18216
rect 34060 18207 34112 18216
rect 34060 18173 34069 18207
rect 34069 18173 34103 18207
rect 34103 18173 34112 18207
rect 34060 18164 34112 18173
rect 34336 18207 34388 18216
rect 34336 18173 34345 18207
rect 34345 18173 34379 18207
rect 34379 18173 34388 18207
rect 34336 18164 34388 18173
rect 18236 18028 18288 18080
rect 19156 18028 19208 18080
rect 25228 18028 25280 18080
rect 27988 18028 28040 18080
rect 28632 18096 28684 18148
rect 29184 18028 29236 18080
rect 31760 18028 31812 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 10600 17867 10652 17876
rect 10600 17833 10609 17867
rect 10609 17833 10643 17867
rect 10643 17833 10652 17867
rect 10600 17824 10652 17833
rect 11060 17824 11112 17876
rect 14280 17867 14332 17876
rect 14280 17833 14289 17867
rect 14289 17833 14323 17867
rect 14323 17833 14332 17867
rect 14280 17824 14332 17833
rect 20168 17824 20220 17876
rect 18696 17756 18748 17808
rect 21824 17824 21876 17876
rect 21916 17824 21968 17876
rect 24584 17867 24636 17876
rect 15844 17688 15896 17740
rect 16212 17731 16264 17740
rect 16212 17697 16221 17731
rect 16221 17697 16255 17731
rect 16255 17697 16264 17731
rect 16212 17688 16264 17697
rect 9772 17620 9824 17672
rect 10600 17663 10652 17672
rect 10600 17629 10609 17663
rect 10609 17629 10643 17663
rect 10643 17629 10652 17663
rect 10600 17620 10652 17629
rect 10784 17663 10836 17672
rect 10784 17629 10793 17663
rect 10793 17629 10827 17663
rect 10827 17629 10836 17663
rect 10784 17620 10836 17629
rect 11244 17663 11296 17672
rect 11244 17629 11253 17663
rect 11253 17629 11287 17663
rect 11287 17629 11296 17663
rect 11244 17620 11296 17629
rect 12164 17620 12216 17672
rect 15016 17620 15068 17672
rect 16948 17552 17000 17604
rect 18052 17620 18104 17672
rect 19524 17663 19576 17672
rect 18328 17552 18380 17604
rect 19524 17629 19533 17663
rect 19533 17629 19567 17663
rect 19567 17629 19576 17663
rect 19524 17620 19576 17629
rect 20812 17663 20864 17672
rect 20812 17629 20821 17663
rect 20821 17629 20855 17663
rect 20855 17629 20864 17663
rect 20812 17620 20864 17629
rect 24584 17833 24593 17867
rect 24593 17833 24627 17867
rect 24627 17833 24636 17867
rect 24584 17824 24636 17833
rect 24768 17867 24820 17876
rect 24768 17833 24777 17867
rect 24777 17833 24811 17867
rect 24811 17833 24820 17867
rect 24768 17824 24820 17833
rect 30104 17824 30156 17876
rect 30380 17824 30432 17876
rect 31392 17867 31444 17876
rect 23756 17756 23808 17808
rect 26792 17756 26844 17808
rect 27252 17731 27304 17740
rect 21456 17620 21508 17672
rect 23296 17663 23348 17672
rect 19340 17552 19392 17604
rect 20444 17552 20496 17604
rect 23296 17629 23305 17663
rect 23305 17629 23339 17663
rect 23339 17629 23348 17663
rect 23296 17620 23348 17629
rect 23388 17663 23440 17672
rect 23388 17629 23397 17663
rect 23397 17629 23431 17663
rect 23431 17629 23440 17663
rect 23388 17620 23440 17629
rect 27252 17697 27261 17731
rect 27261 17697 27295 17731
rect 27295 17697 27304 17731
rect 27252 17688 27304 17697
rect 24676 17620 24728 17672
rect 25504 17620 25556 17672
rect 27160 17620 27212 17672
rect 31392 17833 31401 17867
rect 31401 17833 31435 17867
rect 31435 17833 31444 17867
rect 31392 17824 31444 17833
rect 31208 17756 31260 17808
rect 30840 17663 30892 17672
rect 14924 17527 14976 17536
rect 14924 17493 14933 17527
rect 14933 17493 14967 17527
rect 14967 17493 14976 17527
rect 14924 17484 14976 17493
rect 17868 17527 17920 17536
rect 17868 17493 17877 17527
rect 17877 17493 17911 17527
rect 17911 17493 17920 17527
rect 17868 17484 17920 17493
rect 19064 17484 19116 17536
rect 20168 17484 20220 17536
rect 22560 17527 22612 17536
rect 22560 17493 22569 17527
rect 22569 17493 22603 17527
rect 22603 17493 22612 17527
rect 22560 17484 22612 17493
rect 22652 17484 22704 17536
rect 26424 17552 26476 17604
rect 27804 17484 27856 17536
rect 30840 17629 30849 17663
rect 30849 17629 30883 17663
rect 30883 17629 30892 17663
rect 30840 17620 30892 17629
rect 31484 17663 31536 17672
rect 31484 17629 31493 17663
rect 31493 17629 31527 17663
rect 31527 17629 31536 17663
rect 31484 17620 31536 17629
rect 32956 17688 33008 17740
rect 32404 17663 32456 17672
rect 32404 17629 32413 17663
rect 32413 17629 32447 17663
rect 32447 17629 32456 17663
rect 32404 17620 32456 17629
rect 31852 17552 31904 17604
rect 31024 17484 31076 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 12348 17323 12400 17332
rect 12348 17289 12357 17323
rect 12357 17289 12391 17323
rect 12391 17289 12400 17323
rect 12348 17280 12400 17289
rect 16212 17280 16264 17332
rect 11336 17212 11388 17264
rect 10324 17144 10376 17196
rect 12808 17212 12860 17264
rect 14188 17212 14240 17264
rect 12716 17144 12768 17196
rect 12900 17187 12952 17196
rect 12900 17153 12909 17187
rect 12909 17153 12943 17187
rect 12943 17153 12952 17187
rect 12900 17144 12952 17153
rect 14096 17144 14148 17196
rect 14740 17144 14792 17196
rect 13084 17076 13136 17128
rect 14188 17119 14240 17128
rect 14188 17085 14197 17119
rect 14197 17085 14231 17119
rect 14231 17085 14240 17119
rect 14188 17076 14240 17085
rect 16856 17255 16908 17264
rect 16856 17221 16865 17255
rect 16865 17221 16899 17255
rect 16899 17221 16908 17255
rect 16856 17212 16908 17221
rect 16948 17255 17000 17264
rect 16948 17221 16957 17255
rect 16957 17221 16991 17255
rect 16991 17221 17000 17255
rect 16948 17212 17000 17221
rect 17132 17212 17184 17264
rect 18328 17212 18380 17264
rect 17040 17187 17092 17196
rect 17040 17153 17049 17187
rect 17049 17153 17083 17187
rect 17083 17153 17092 17187
rect 17040 17144 17092 17153
rect 19156 17144 19208 17196
rect 22744 17212 22796 17264
rect 17040 17008 17092 17060
rect 20168 17144 20220 17196
rect 19524 17076 19576 17128
rect 20904 17144 20956 17196
rect 22100 17187 22152 17196
rect 22100 17153 22109 17187
rect 22109 17153 22143 17187
rect 22143 17153 22152 17187
rect 22100 17144 22152 17153
rect 23756 17187 23808 17196
rect 23756 17153 23765 17187
rect 23765 17153 23799 17187
rect 23799 17153 23808 17187
rect 23756 17144 23808 17153
rect 25228 17187 25280 17196
rect 25228 17153 25237 17187
rect 25237 17153 25271 17187
rect 25271 17153 25280 17187
rect 25228 17144 25280 17153
rect 21456 17076 21508 17128
rect 12624 16940 12676 16992
rect 17224 16983 17276 16992
rect 17224 16949 17233 16983
rect 17233 16949 17267 16983
rect 17267 16949 17276 16983
rect 17224 16940 17276 16949
rect 18144 16940 18196 16992
rect 19432 16940 19484 16992
rect 20260 16940 20312 16992
rect 22836 16983 22888 16992
rect 22836 16949 22845 16983
rect 22845 16949 22879 16983
rect 22879 16949 22888 16983
rect 22836 16940 22888 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 10600 16736 10652 16788
rect 12808 16779 12860 16788
rect 12808 16745 12817 16779
rect 12817 16745 12851 16779
rect 12851 16745 12860 16779
rect 12808 16736 12860 16745
rect 14188 16736 14240 16788
rect 9404 16600 9456 16652
rect 12716 16668 12768 16720
rect 14740 16711 14792 16720
rect 14740 16677 14749 16711
rect 14749 16677 14783 16711
rect 14783 16677 14792 16711
rect 14740 16668 14792 16677
rect 13084 16600 13136 16652
rect 20076 16736 20128 16788
rect 16948 16668 17000 16720
rect 18236 16668 18288 16720
rect 20996 16668 21048 16720
rect 12624 16575 12676 16584
rect 12624 16541 12633 16575
rect 12633 16541 12667 16575
rect 12667 16541 12676 16575
rect 12900 16575 12952 16584
rect 12624 16532 12676 16541
rect 12900 16541 12909 16575
rect 12909 16541 12943 16575
rect 12943 16541 12952 16575
rect 12900 16532 12952 16541
rect 13544 16575 13596 16584
rect 13544 16541 13553 16575
rect 13553 16541 13587 16575
rect 13587 16541 13596 16575
rect 13544 16532 13596 16541
rect 14096 16575 14148 16584
rect 14096 16541 14105 16575
rect 14105 16541 14139 16575
rect 14139 16541 14148 16575
rect 14096 16532 14148 16541
rect 14924 16575 14976 16584
rect 14924 16541 14933 16575
rect 14933 16541 14967 16575
rect 14967 16541 14976 16575
rect 14924 16532 14976 16541
rect 17224 16532 17276 16584
rect 17868 16575 17920 16584
rect 17868 16541 17877 16575
rect 17877 16541 17911 16575
rect 17911 16541 17920 16575
rect 17868 16532 17920 16541
rect 18696 16575 18748 16584
rect 18696 16541 18705 16575
rect 18705 16541 18739 16575
rect 18739 16541 18748 16575
rect 18696 16532 18748 16541
rect 19340 16575 19392 16584
rect 19340 16541 19349 16575
rect 19349 16541 19383 16575
rect 19383 16541 19392 16575
rect 19340 16532 19392 16541
rect 21456 16575 21508 16584
rect 9588 16464 9640 16516
rect 19156 16464 19208 16516
rect 21456 16541 21465 16575
rect 21465 16541 21499 16575
rect 21499 16541 21508 16575
rect 21456 16532 21508 16541
rect 23020 16532 23072 16584
rect 23756 16532 23808 16584
rect 25412 16575 25464 16584
rect 25412 16541 25421 16575
rect 25421 16541 25455 16575
rect 25455 16541 25464 16575
rect 25412 16532 25464 16541
rect 11796 16396 11848 16448
rect 13360 16439 13412 16448
rect 13360 16405 13369 16439
rect 13369 16405 13403 16439
rect 13403 16405 13412 16439
rect 13360 16396 13412 16405
rect 18696 16396 18748 16448
rect 22468 16439 22520 16448
rect 22468 16405 22477 16439
rect 22477 16405 22511 16439
rect 22511 16405 22520 16439
rect 22468 16396 22520 16405
rect 23204 16439 23256 16448
rect 23204 16405 23213 16439
rect 23213 16405 23247 16439
rect 23247 16405 23256 16439
rect 23204 16396 23256 16405
rect 23480 16396 23532 16448
rect 24400 16396 24452 16448
rect 25688 16396 25740 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 12624 16192 12676 16244
rect 14096 16192 14148 16244
rect 16488 16235 16540 16244
rect 16488 16201 16497 16235
rect 16497 16201 16531 16235
rect 16531 16201 16540 16235
rect 16488 16192 16540 16201
rect 19340 16192 19392 16244
rect 22560 16192 22612 16244
rect 9404 16124 9456 16176
rect 13360 16124 13412 16176
rect 8300 16056 8352 16108
rect 8576 16099 8628 16108
rect 8576 16065 8585 16099
rect 8585 16065 8619 16099
rect 8619 16065 8628 16099
rect 8576 16056 8628 16065
rect 8852 16099 8904 16108
rect 8852 16065 8886 16099
rect 8886 16065 8904 16099
rect 8852 16056 8904 16065
rect 13176 16056 13228 16108
rect 14188 16056 14240 16108
rect 12256 15988 12308 16040
rect 11796 15963 11848 15972
rect 11796 15929 11805 15963
rect 11805 15929 11839 15963
rect 11839 15929 11848 15963
rect 11796 15920 11848 15929
rect 18696 16099 18748 16108
rect 18696 16065 18705 16099
rect 18705 16065 18739 16099
rect 18739 16065 18748 16099
rect 18696 16056 18748 16065
rect 19340 16056 19392 16108
rect 20260 16099 20312 16108
rect 20260 16065 20269 16099
rect 20269 16065 20303 16099
rect 20303 16065 20312 16099
rect 20260 16056 20312 16065
rect 25044 16192 25096 16244
rect 25412 16192 25464 16244
rect 23204 16124 23256 16176
rect 23480 16056 23532 16108
rect 25504 16056 25556 16108
rect 25688 16056 25740 16108
rect 26056 16099 26108 16108
rect 26056 16065 26065 16099
rect 26065 16065 26099 16099
rect 26099 16065 26108 16099
rect 26056 16056 26108 16065
rect 18052 15988 18104 16040
rect 19156 15988 19208 16040
rect 22928 16031 22980 16040
rect 22928 15997 22937 16031
rect 22937 15997 22971 16031
rect 22971 15997 22980 16031
rect 22928 15988 22980 15997
rect 16396 15920 16448 15972
rect 18880 15920 18932 15972
rect 7748 15895 7800 15904
rect 7748 15861 7757 15895
rect 7757 15861 7791 15895
rect 7791 15861 7800 15895
rect 7748 15852 7800 15861
rect 9956 15895 10008 15904
rect 9956 15861 9965 15895
rect 9965 15861 9999 15895
rect 9999 15861 10008 15895
rect 9956 15852 10008 15861
rect 17592 15895 17644 15904
rect 17592 15861 17601 15895
rect 17601 15861 17635 15895
rect 17635 15861 17644 15895
rect 17592 15852 17644 15861
rect 22100 15852 22152 15904
rect 23572 15852 23624 15904
rect 26240 15852 26292 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 8576 15648 8628 15700
rect 8852 15648 8904 15700
rect 9588 15691 9640 15700
rect 9588 15657 9597 15691
rect 9597 15657 9631 15691
rect 9631 15657 9640 15691
rect 9588 15648 9640 15657
rect 12900 15648 12952 15700
rect 13544 15648 13596 15700
rect 12256 15580 12308 15632
rect 18236 15648 18288 15700
rect 7012 15555 7064 15564
rect 7012 15521 7021 15555
rect 7021 15521 7055 15555
rect 7055 15521 7064 15555
rect 7012 15512 7064 15521
rect 9956 15555 10008 15564
rect 9956 15521 9965 15555
rect 9965 15521 9999 15555
rect 9999 15521 10008 15555
rect 9956 15512 10008 15521
rect 7748 15444 7800 15496
rect 9128 15487 9180 15496
rect 9128 15453 9137 15487
rect 9137 15453 9171 15487
rect 9171 15453 9180 15487
rect 9128 15444 9180 15453
rect 9772 15487 9824 15496
rect 9772 15453 9781 15487
rect 9781 15453 9815 15487
rect 9815 15453 9824 15487
rect 9772 15444 9824 15453
rect 9864 15487 9916 15496
rect 9864 15453 9873 15487
rect 9873 15453 9907 15487
rect 9907 15453 9916 15487
rect 10876 15487 10928 15496
rect 9864 15444 9916 15453
rect 10876 15453 10885 15487
rect 10885 15453 10919 15487
rect 10919 15453 10928 15487
rect 10876 15444 10928 15453
rect 11796 15512 11848 15564
rect 19156 15580 19208 15632
rect 21456 15648 21508 15700
rect 23756 15691 23808 15700
rect 23756 15657 23765 15691
rect 23765 15657 23799 15691
rect 23799 15657 23808 15691
rect 23756 15648 23808 15657
rect 25044 15691 25096 15700
rect 25044 15657 25053 15691
rect 25053 15657 25087 15691
rect 25087 15657 25096 15691
rect 25044 15648 25096 15657
rect 26056 15648 26108 15700
rect 22468 15512 22520 15564
rect 10140 15376 10192 15428
rect 11336 15444 11388 15496
rect 13452 15444 13504 15496
rect 15016 15444 15068 15496
rect 17960 15487 18012 15496
rect 17960 15453 17969 15487
rect 17969 15453 18003 15487
rect 18003 15453 18012 15487
rect 17960 15444 18012 15453
rect 19432 15444 19484 15496
rect 21088 15444 21140 15496
rect 22376 15444 22428 15496
rect 22928 15512 22980 15564
rect 23572 15487 23624 15496
rect 16672 15376 16724 15428
rect 22744 15376 22796 15428
rect 23572 15453 23581 15487
rect 23581 15453 23615 15487
rect 23615 15453 23624 15487
rect 23572 15444 23624 15453
rect 8392 15351 8444 15360
rect 8392 15317 8401 15351
rect 8401 15317 8435 15351
rect 8435 15317 8444 15351
rect 8392 15308 8444 15317
rect 9588 15308 9640 15360
rect 15200 15308 15252 15360
rect 18420 15308 18472 15360
rect 20260 15351 20312 15360
rect 20260 15317 20269 15351
rect 20269 15317 20303 15351
rect 20303 15317 20312 15351
rect 20260 15308 20312 15317
rect 20812 15308 20864 15360
rect 22468 15308 22520 15360
rect 23940 15308 23992 15360
rect 25320 15308 25372 15360
rect 25504 15444 25556 15496
rect 25504 15308 25556 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 8300 15147 8352 15156
rect 8300 15113 8309 15147
rect 8309 15113 8343 15147
rect 8343 15113 8352 15147
rect 8300 15104 8352 15113
rect 9128 15147 9180 15156
rect 9128 15113 9137 15147
rect 9137 15113 9171 15147
rect 9171 15113 9180 15147
rect 9128 15104 9180 15113
rect 16672 15147 16724 15156
rect 8392 15036 8444 15088
rect 9956 15036 10008 15088
rect 8024 14900 8076 14952
rect 6920 14764 6972 14816
rect 9404 14968 9456 15020
rect 9864 15011 9916 15020
rect 9864 14977 9898 15011
rect 9898 14977 9916 15011
rect 9864 14968 9916 14977
rect 10232 14968 10284 15020
rect 12440 15036 12492 15088
rect 16672 15113 16681 15147
rect 16681 15113 16715 15147
rect 16715 15113 16724 15147
rect 16672 15104 16724 15113
rect 23940 15147 23992 15156
rect 18236 15036 18288 15088
rect 20996 15079 21048 15088
rect 20996 15045 21005 15079
rect 21005 15045 21039 15079
rect 21039 15045 21048 15079
rect 20996 15036 21048 15045
rect 23940 15113 23949 15147
rect 23949 15113 23983 15147
rect 23983 15113 23992 15147
rect 23940 15104 23992 15113
rect 25688 15104 25740 15156
rect 12716 15011 12768 15020
rect 10600 14900 10652 14952
rect 12716 14977 12725 15011
rect 12725 14977 12759 15011
rect 12759 14977 12768 15011
rect 12716 14968 12768 14977
rect 15200 14968 15252 15020
rect 17592 14968 17644 15020
rect 19984 14968 20036 15020
rect 20352 14968 20404 15020
rect 13176 14943 13228 14952
rect 13176 14909 13185 14943
rect 13185 14909 13219 14943
rect 13219 14909 13228 14943
rect 13176 14900 13228 14909
rect 19156 14900 19208 14952
rect 23112 14968 23164 15020
rect 22376 14900 22428 14952
rect 10968 14807 11020 14816
rect 10968 14773 10977 14807
rect 10977 14773 11011 14807
rect 11011 14773 11020 14807
rect 10968 14764 11020 14773
rect 11704 14764 11756 14816
rect 14556 14807 14608 14816
rect 14556 14773 14565 14807
rect 14565 14773 14599 14807
rect 14599 14773 14608 14807
rect 14556 14764 14608 14773
rect 18972 14764 19024 14816
rect 20444 14807 20496 14816
rect 20444 14773 20453 14807
rect 20453 14773 20487 14807
rect 20487 14773 20496 14807
rect 20444 14764 20496 14773
rect 21088 14807 21140 14816
rect 21088 14773 21097 14807
rect 21097 14773 21131 14807
rect 21131 14773 21140 14807
rect 21088 14764 21140 14773
rect 21364 14764 21416 14816
rect 25320 14968 25372 15020
rect 24308 14900 24360 14952
rect 25228 14900 25280 14952
rect 25412 14943 25464 14952
rect 25412 14909 25421 14943
rect 25421 14909 25455 14943
rect 25455 14909 25464 14943
rect 25412 14900 25464 14909
rect 25044 14832 25096 14884
rect 26056 14968 26108 15020
rect 25964 14764 26016 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 7012 14560 7064 14612
rect 9588 14560 9640 14612
rect 9772 14560 9824 14612
rect 10600 14603 10652 14612
rect 10600 14569 10609 14603
rect 10609 14569 10643 14603
rect 10643 14569 10652 14603
rect 10600 14560 10652 14569
rect 10876 14560 10928 14612
rect 13084 14603 13136 14612
rect 13084 14569 13093 14603
rect 13093 14569 13127 14603
rect 13127 14569 13136 14603
rect 13084 14560 13136 14569
rect 15384 14560 15436 14612
rect 16396 14603 16448 14612
rect 16396 14569 16405 14603
rect 16405 14569 16439 14603
rect 16439 14569 16448 14603
rect 16396 14560 16448 14569
rect 18880 14560 18932 14612
rect 23112 14603 23164 14612
rect 23112 14569 23121 14603
rect 23121 14569 23155 14603
rect 23155 14569 23164 14603
rect 23112 14560 23164 14569
rect 23940 14560 23992 14612
rect 9956 14424 10008 14476
rect 11060 14424 11112 14476
rect 6920 14356 6972 14408
rect 10968 14356 11020 14408
rect 14556 14424 14608 14476
rect 9588 14288 9640 14340
rect 11520 14288 11572 14340
rect 12440 14356 12492 14408
rect 12900 14356 12952 14408
rect 15016 14399 15068 14408
rect 15016 14365 15048 14399
rect 15048 14365 15068 14399
rect 15016 14356 15068 14365
rect 15568 14356 15620 14408
rect 17316 14399 17368 14408
rect 17316 14365 17325 14399
rect 17325 14365 17359 14399
rect 17359 14365 17368 14399
rect 17316 14356 17368 14365
rect 19432 14399 19484 14408
rect 19432 14365 19441 14399
rect 19441 14365 19475 14399
rect 19475 14365 19484 14399
rect 19432 14356 19484 14365
rect 21364 14356 21416 14408
rect 22284 14424 22336 14476
rect 22468 14424 22520 14476
rect 22744 14399 22796 14408
rect 13176 14288 13228 14340
rect 15292 14331 15344 14340
rect 15292 14297 15326 14331
rect 15326 14297 15344 14331
rect 15292 14288 15344 14297
rect 8300 14220 8352 14272
rect 9956 14220 10008 14272
rect 16120 14220 16172 14272
rect 19984 14288 20036 14340
rect 19340 14220 19392 14272
rect 21824 14288 21876 14340
rect 22744 14365 22753 14399
rect 22753 14365 22787 14399
rect 22787 14365 22796 14399
rect 22744 14356 22796 14365
rect 24676 14356 24728 14408
rect 25044 14467 25096 14476
rect 25044 14433 25053 14467
rect 25053 14433 25087 14467
rect 25087 14433 25096 14467
rect 25044 14424 25096 14433
rect 25688 14424 25740 14476
rect 26240 14399 26292 14408
rect 26240 14365 26274 14399
rect 26274 14365 26292 14399
rect 26240 14356 26292 14365
rect 21456 14263 21508 14272
rect 21456 14229 21465 14263
rect 21465 14229 21499 14263
rect 21499 14229 21508 14263
rect 24308 14288 24360 14340
rect 22284 14263 22336 14272
rect 21456 14220 21508 14229
rect 22284 14229 22293 14263
rect 22293 14229 22327 14263
rect 22327 14229 22336 14263
rect 22284 14220 22336 14229
rect 24124 14220 24176 14272
rect 25228 14288 25280 14340
rect 25412 14220 25464 14272
rect 37740 14220 37792 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 9956 14059 10008 14068
rect 9956 14025 9965 14059
rect 9965 14025 9999 14059
rect 9999 14025 10008 14059
rect 9956 14016 10008 14025
rect 10232 14016 10284 14068
rect 12716 14016 12768 14068
rect 18972 14059 19024 14068
rect 8300 13948 8352 14000
rect 9772 13991 9824 14000
rect 9772 13957 9781 13991
rect 9781 13957 9815 13991
rect 9815 13957 9824 13991
rect 9772 13948 9824 13957
rect 8024 13880 8076 13932
rect 8760 13923 8812 13932
rect 8484 13812 8536 13864
rect 8760 13889 8769 13923
rect 8769 13889 8803 13923
rect 8803 13889 8812 13923
rect 8760 13880 8812 13889
rect 9588 13923 9640 13932
rect 9588 13889 9597 13923
rect 9597 13889 9631 13923
rect 9631 13889 9640 13923
rect 9588 13880 9640 13889
rect 9680 13923 9732 13932
rect 9680 13889 9689 13923
rect 9689 13889 9723 13923
rect 9723 13889 9732 13923
rect 11612 13948 11664 14000
rect 15384 13948 15436 14000
rect 9680 13880 9732 13889
rect 11704 13923 11756 13932
rect 11704 13889 11713 13923
rect 11713 13889 11747 13923
rect 11747 13889 11756 13923
rect 11704 13880 11756 13889
rect 12624 13880 12676 13932
rect 12900 13880 12952 13932
rect 13452 13923 13504 13932
rect 13452 13889 13461 13923
rect 13461 13889 13495 13923
rect 13495 13889 13504 13923
rect 13452 13880 13504 13889
rect 15108 13923 15160 13932
rect 15108 13889 15117 13923
rect 15117 13889 15151 13923
rect 15151 13889 15160 13923
rect 15108 13880 15160 13889
rect 18972 14025 18981 14059
rect 18981 14025 19015 14059
rect 19015 14025 19024 14059
rect 18972 14016 19024 14025
rect 19984 14016 20036 14068
rect 20352 14059 20404 14068
rect 20352 14025 20361 14059
rect 20361 14025 20395 14059
rect 20395 14025 20404 14059
rect 20352 14016 20404 14025
rect 21456 14016 21508 14068
rect 22192 14016 22244 14068
rect 22836 14016 22888 14068
rect 26516 14016 26568 14068
rect 18880 13991 18932 14000
rect 18880 13957 18889 13991
rect 18889 13957 18923 13991
rect 18923 13957 18932 13991
rect 18880 13948 18932 13957
rect 20812 13991 20864 14000
rect 20812 13957 20821 13991
rect 20821 13957 20855 13991
rect 20855 13957 20864 13991
rect 20812 13948 20864 13957
rect 24860 13948 24912 14000
rect 25504 13948 25556 14000
rect 16120 13923 16172 13932
rect 9128 13812 9180 13864
rect 13268 13855 13320 13864
rect 13268 13821 13277 13855
rect 13277 13821 13311 13855
rect 13311 13821 13320 13855
rect 13268 13812 13320 13821
rect 15384 13812 15436 13864
rect 16120 13889 16129 13923
rect 16129 13889 16163 13923
rect 16163 13889 16172 13923
rect 16120 13880 16172 13889
rect 17132 13880 17184 13932
rect 18052 13880 18104 13932
rect 20444 13880 20496 13932
rect 22376 13923 22428 13932
rect 22376 13889 22385 13923
rect 22385 13889 22419 13923
rect 22419 13889 22428 13923
rect 22376 13880 22428 13889
rect 24124 13923 24176 13932
rect 24124 13889 24133 13923
rect 24133 13889 24167 13923
rect 24167 13889 24176 13923
rect 24124 13880 24176 13889
rect 24952 13880 25004 13932
rect 25044 13880 25096 13932
rect 26056 13991 26108 14000
rect 26056 13957 26081 13991
rect 26081 13957 26108 13991
rect 26056 13948 26108 13957
rect 11796 13744 11848 13796
rect 3792 13676 3844 13728
rect 10232 13676 10284 13728
rect 14924 13676 14976 13728
rect 17960 13744 18012 13796
rect 18604 13744 18656 13796
rect 21088 13812 21140 13864
rect 22468 13812 22520 13864
rect 23756 13855 23808 13864
rect 23756 13821 23765 13855
rect 23765 13821 23799 13855
rect 23799 13821 23808 13855
rect 23756 13812 23808 13821
rect 24216 13855 24268 13864
rect 24216 13821 24225 13855
rect 24225 13821 24259 13855
rect 24259 13821 24268 13855
rect 24216 13812 24268 13821
rect 25228 13812 25280 13864
rect 26792 13744 26844 13796
rect 27620 13787 27672 13796
rect 27620 13753 27629 13787
rect 27629 13753 27663 13787
rect 27663 13753 27672 13787
rect 27620 13744 27672 13753
rect 15752 13676 15804 13728
rect 18052 13676 18104 13728
rect 23664 13676 23716 13728
rect 25228 13719 25280 13728
rect 25228 13685 25237 13719
rect 25237 13685 25271 13719
rect 25271 13685 25280 13719
rect 25228 13676 25280 13685
rect 25964 13676 26016 13728
rect 26148 13676 26200 13728
rect 26424 13676 26476 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 8760 13472 8812 13524
rect 9588 13472 9640 13524
rect 10140 13515 10192 13524
rect 10140 13481 10149 13515
rect 10149 13481 10183 13515
rect 10183 13481 10192 13515
rect 10140 13472 10192 13481
rect 10232 13472 10284 13524
rect 7012 13379 7064 13388
rect 7012 13345 7021 13379
rect 7021 13345 7055 13379
rect 7055 13345 7064 13379
rect 7012 13336 7064 13345
rect 9680 13336 9732 13388
rect 8484 13268 8536 13320
rect 15292 13404 15344 13456
rect 19432 13404 19484 13456
rect 24952 13404 25004 13456
rect 25596 13404 25648 13456
rect 26148 13404 26200 13456
rect 11612 13311 11664 13320
rect 11612 13277 11621 13311
rect 11621 13277 11655 13311
rect 11655 13277 11664 13311
rect 11612 13268 11664 13277
rect 14556 13336 14608 13388
rect 15108 13336 15160 13388
rect 17960 13336 18012 13388
rect 18144 13336 18196 13388
rect 19248 13379 19300 13388
rect 19248 13345 19257 13379
rect 19257 13345 19291 13379
rect 19291 13345 19300 13379
rect 19248 13336 19300 13345
rect 25044 13379 25096 13388
rect 9772 13200 9824 13252
rect 10968 13200 11020 13252
rect 11796 13243 11848 13252
rect 11796 13209 11805 13243
rect 11805 13209 11839 13243
rect 11839 13209 11848 13243
rect 11796 13200 11848 13209
rect 13452 13268 13504 13320
rect 14556 13200 14608 13252
rect 12532 13175 12584 13184
rect 12532 13141 12541 13175
rect 12541 13141 12575 13175
rect 12575 13141 12584 13175
rect 12532 13132 12584 13141
rect 14740 13311 14792 13320
rect 14740 13277 14749 13311
rect 14749 13277 14783 13311
rect 14783 13277 14792 13311
rect 14924 13311 14976 13320
rect 14740 13268 14792 13277
rect 14924 13277 14926 13311
rect 14926 13277 14960 13311
rect 14960 13277 14976 13311
rect 14924 13268 14976 13277
rect 15752 13311 15804 13320
rect 15752 13277 15786 13311
rect 15786 13277 15804 13311
rect 15752 13268 15804 13277
rect 18052 13311 18104 13320
rect 18052 13277 18061 13311
rect 18061 13277 18095 13311
rect 18095 13277 18104 13311
rect 18052 13268 18104 13277
rect 19432 13311 19484 13320
rect 19432 13277 19441 13311
rect 19441 13277 19475 13311
rect 19475 13277 19484 13311
rect 19432 13268 19484 13277
rect 21088 13268 21140 13320
rect 21364 13268 21416 13320
rect 22284 13268 22336 13320
rect 25044 13345 25053 13379
rect 25053 13345 25087 13379
rect 25087 13345 25096 13379
rect 25044 13336 25096 13345
rect 24768 13268 24820 13320
rect 26332 13336 26384 13388
rect 16948 13200 17000 13252
rect 15108 13132 15160 13184
rect 15660 13132 15712 13184
rect 17960 13132 18012 13184
rect 19248 13132 19300 13184
rect 25688 13200 25740 13252
rect 26148 13200 26200 13252
rect 26332 13243 26384 13252
rect 26332 13209 26341 13243
rect 26341 13209 26375 13243
rect 26375 13209 26384 13243
rect 26332 13200 26384 13209
rect 26976 13268 27028 13320
rect 27160 13200 27212 13252
rect 22376 13132 22428 13184
rect 23388 13132 23440 13184
rect 24124 13132 24176 13184
rect 24952 13132 25004 13184
rect 25504 13132 25556 13184
rect 25780 13132 25832 13184
rect 27620 13132 27672 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 1492 12860 1544 12912
rect 12532 12860 12584 12912
rect 15476 12928 15528 12980
rect 20260 12928 20312 12980
rect 22100 12928 22152 12980
rect 26332 12928 26384 12980
rect 7012 12792 7064 12844
rect 8116 12792 8168 12844
rect 8852 12792 8904 12844
rect 9956 12835 10008 12844
rect 9956 12801 9965 12835
rect 9965 12801 9999 12835
rect 9999 12801 10008 12835
rect 9956 12792 10008 12801
rect 9680 12724 9732 12776
rect 11612 12792 11664 12844
rect 12348 12792 12400 12844
rect 14740 12792 14792 12844
rect 15476 12835 15528 12844
rect 15476 12801 15485 12835
rect 15485 12801 15519 12835
rect 15519 12801 15528 12835
rect 15476 12792 15528 12801
rect 11520 12767 11572 12776
rect 11520 12733 11529 12767
rect 11529 12733 11563 12767
rect 11563 12733 11572 12767
rect 11520 12724 11572 12733
rect 13176 12724 13228 12776
rect 14556 12724 14608 12776
rect 15660 12724 15712 12776
rect 11060 12656 11112 12708
rect 9680 12588 9732 12640
rect 13268 12588 13320 12640
rect 14556 12588 14608 12640
rect 14740 12631 14792 12640
rect 14740 12597 14749 12631
rect 14749 12597 14783 12631
rect 14783 12597 14792 12631
rect 14740 12588 14792 12597
rect 15568 12588 15620 12640
rect 18144 12860 18196 12912
rect 20904 12860 20956 12912
rect 16948 12792 17000 12844
rect 20628 12792 20680 12844
rect 16764 12724 16816 12776
rect 17316 12767 17368 12776
rect 17316 12733 17325 12767
rect 17325 12733 17359 12767
rect 17359 12733 17368 12767
rect 17316 12724 17368 12733
rect 18604 12724 18656 12776
rect 22192 12835 22244 12844
rect 22192 12801 22201 12835
rect 22201 12801 22235 12835
rect 22235 12801 22244 12835
rect 22192 12792 22244 12801
rect 23664 12835 23716 12844
rect 23664 12801 23673 12835
rect 23673 12801 23707 12835
rect 23707 12801 23716 12835
rect 23664 12792 23716 12801
rect 24124 12835 24176 12844
rect 24124 12801 24133 12835
rect 24133 12801 24167 12835
rect 24167 12801 24176 12835
rect 24124 12792 24176 12801
rect 24952 12835 25004 12844
rect 24952 12801 24961 12835
rect 24961 12801 24995 12835
rect 24995 12801 25004 12835
rect 24952 12792 25004 12801
rect 26240 12860 26292 12912
rect 24216 12724 24268 12776
rect 24768 12724 24820 12776
rect 24584 12656 24636 12708
rect 25780 12724 25832 12776
rect 26424 12835 26476 12844
rect 26424 12801 26433 12835
rect 26433 12801 26467 12835
rect 26467 12801 26476 12835
rect 26976 12835 27028 12844
rect 26424 12792 26476 12801
rect 26976 12801 26985 12835
rect 26985 12801 27019 12835
rect 27019 12801 27028 12835
rect 26976 12792 27028 12801
rect 27160 12835 27212 12844
rect 27160 12801 27169 12835
rect 27169 12801 27203 12835
rect 27203 12801 27212 12835
rect 27160 12792 27212 12801
rect 26516 12724 26568 12776
rect 26792 12724 26844 12776
rect 27620 12860 27672 12912
rect 28172 12835 28224 12844
rect 18696 12631 18748 12640
rect 18696 12597 18705 12631
rect 18705 12597 18739 12631
rect 18739 12597 18748 12631
rect 18696 12588 18748 12597
rect 19340 12588 19392 12640
rect 21824 12631 21876 12640
rect 21824 12597 21833 12631
rect 21833 12597 21867 12631
rect 21867 12597 21876 12631
rect 21824 12588 21876 12597
rect 24768 12588 24820 12640
rect 26240 12656 26292 12708
rect 28172 12801 28181 12835
rect 28181 12801 28215 12835
rect 28215 12801 28224 12835
rect 28172 12792 28224 12801
rect 37832 12835 37884 12844
rect 37832 12801 37841 12835
rect 37841 12801 37875 12835
rect 37875 12801 37884 12835
rect 37832 12792 37884 12801
rect 38200 12656 38252 12708
rect 38016 12631 38068 12640
rect 38016 12597 38025 12631
rect 38025 12597 38059 12631
rect 38059 12597 38068 12631
rect 38016 12588 38068 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 8852 12384 8904 12436
rect 10968 12427 11020 12436
rect 10968 12393 10977 12427
rect 10977 12393 11011 12427
rect 11011 12393 11020 12427
rect 10968 12384 11020 12393
rect 12440 12384 12492 12436
rect 14740 12384 14792 12436
rect 15292 12427 15344 12436
rect 15292 12393 15301 12427
rect 15301 12393 15335 12427
rect 15335 12393 15344 12427
rect 15292 12384 15344 12393
rect 17224 12427 17276 12436
rect 17224 12393 17233 12427
rect 17233 12393 17267 12427
rect 17267 12393 17276 12427
rect 17224 12384 17276 12393
rect 19432 12384 19484 12436
rect 20628 12427 20680 12436
rect 20628 12393 20637 12427
rect 20637 12393 20671 12427
rect 20671 12393 20680 12427
rect 20628 12384 20680 12393
rect 27620 12384 27672 12436
rect 28172 12384 28224 12436
rect 11612 12316 11664 12368
rect 8116 12248 8168 12300
rect 11796 12248 11848 12300
rect 12256 12291 12308 12300
rect 12256 12257 12265 12291
rect 12265 12257 12299 12291
rect 12299 12257 12308 12291
rect 12256 12248 12308 12257
rect 15200 12316 15252 12368
rect 9128 12223 9180 12232
rect 9128 12189 9137 12223
rect 9137 12189 9171 12223
rect 9171 12189 9180 12223
rect 9128 12180 9180 12189
rect 14740 12248 14792 12300
rect 18420 12291 18472 12300
rect 18420 12257 18429 12291
rect 18429 12257 18463 12291
rect 18463 12257 18472 12291
rect 18420 12248 18472 12257
rect 18604 12291 18656 12300
rect 18604 12257 18613 12291
rect 18613 12257 18647 12291
rect 18647 12257 18656 12291
rect 18604 12248 18656 12257
rect 18696 12248 18748 12300
rect 9496 12112 9548 12164
rect 11244 12112 11296 12164
rect 13452 12180 13504 12232
rect 14648 12180 14700 12232
rect 14556 12112 14608 12164
rect 15476 12112 15528 12164
rect 16488 12112 16540 12164
rect 17316 12112 17368 12164
rect 14280 12044 14332 12096
rect 14740 12044 14792 12096
rect 21364 12180 21416 12232
rect 23388 12291 23440 12300
rect 23388 12257 23397 12291
rect 23397 12257 23431 12291
rect 23431 12257 23440 12291
rect 23388 12248 23440 12257
rect 25412 12316 25464 12368
rect 26240 12316 26292 12368
rect 23756 12248 23808 12300
rect 24584 12248 24636 12300
rect 22192 12180 22244 12232
rect 23572 12180 23624 12232
rect 25872 12180 25924 12232
rect 26424 12180 26476 12232
rect 26608 12223 26660 12232
rect 26608 12189 26617 12223
rect 26617 12189 26651 12223
rect 26651 12189 26660 12223
rect 27068 12223 27120 12232
rect 26608 12180 26660 12189
rect 27068 12189 27077 12223
rect 27077 12189 27111 12223
rect 27111 12189 27120 12223
rect 27068 12180 27120 12189
rect 20720 12044 20772 12096
rect 20996 12044 21048 12096
rect 21732 12087 21784 12096
rect 21732 12053 21741 12087
rect 21741 12053 21775 12087
rect 21775 12053 21784 12087
rect 21732 12044 21784 12053
rect 37832 12112 37884 12164
rect 22744 12044 22796 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 9496 11883 9548 11892
rect 9496 11849 9505 11883
rect 9505 11849 9539 11883
rect 9539 11849 9548 11883
rect 9496 11840 9548 11849
rect 21364 11840 21416 11892
rect 27160 11840 27212 11892
rect 8668 11747 8720 11756
rect 8668 11713 8677 11747
rect 8677 11713 8711 11747
rect 8711 11713 8720 11747
rect 8668 11704 8720 11713
rect 9680 11747 9732 11756
rect 9680 11713 9689 11747
rect 9689 11713 9723 11747
rect 9723 11713 9732 11747
rect 9680 11704 9732 11713
rect 8208 11636 8260 11688
rect 10324 11636 10376 11688
rect 12624 11704 12676 11756
rect 12900 11704 12952 11756
rect 13452 11704 13504 11756
rect 14280 11747 14332 11756
rect 14280 11713 14289 11747
rect 14289 11713 14323 11747
rect 14323 11713 14332 11747
rect 14280 11704 14332 11713
rect 14832 11704 14884 11756
rect 16488 11704 16540 11756
rect 19340 11747 19392 11756
rect 19340 11713 19349 11747
rect 19349 11713 19383 11747
rect 19383 11713 19392 11747
rect 19340 11704 19392 11713
rect 21824 11772 21876 11824
rect 21732 11704 21784 11756
rect 23480 11704 23532 11756
rect 14648 11636 14700 11688
rect 16120 11636 16172 11688
rect 19248 11636 19300 11688
rect 22744 11679 22796 11688
rect 22744 11645 22753 11679
rect 22753 11645 22787 11679
rect 22787 11645 22796 11679
rect 22744 11636 22796 11645
rect 23572 11636 23624 11688
rect 24216 11636 24268 11688
rect 26056 11704 26108 11756
rect 26424 11704 26476 11756
rect 27068 11704 27120 11756
rect 27620 11747 27672 11756
rect 27620 11713 27629 11747
rect 27629 11713 27663 11747
rect 27663 11713 27672 11747
rect 27620 11704 27672 11713
rect 25964 11679 26016 11688
rect 25964 11645 25973 11679
rect 25973 11645 26007 11679
rect 26007 11645 26016 11679
rect 25964 11636 26016 11645
rect 26240 11636 26292 11688
rect 21916 11568 21968 11620
rect 26792 11568 26844 11620
rect 9036 11500 9088 11552
rect 11336 11500 11388 11552
rect 12164 11500 12216 11552
rect 15476 11500 15528 11552
rect 20812 11543 20864 11552
rect 20812 11509 20821 11543
rect 20821 11509 20855 11543
rect 20855 11509 20864 11543
rect 20812 11500 20864 11509
rect 24124 11500 24176 11552
rect 24216 11500 24268 11552
rect 25320 11500 25372 11552
rect 26148 11500 26200 11552
rect 26332 11500 26384 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 12256 11296 12308 11348
rect 14740 11339 14792 11348
rect 14740 11305 14749 11339
rect 14749 11305 14783 11339
rect 14783 11305 14792 11339
rect 14740 11296 14792 11305
rect 18144 11271 18196 11280
rect 12900 11160 12952 11212
rect 16672 11160 16724 11212
rect 18144 11237 18153 11271
rect 18153 11237 18187 11271
rect 18187 11237 18196 11271
rect 18144 11228 18196 11237
rect 18512 11228 18564 11280
rect 19340 11228 19392 11280
rect 22192 11228 22244 11280
rect 24676 11228 24728 11280
rect 26424 11228 26476 11280
rect 20720 11203 20772 11212
rect 8116 11092 8168 11144
rect 7564 11024 7616 11076
rect 9036 11092 9088 11144
rect 10232 11092 10284 11144
rect 10876 11092 10928 11144
rect 1584 10999 1636 11008
rect 1584 10965 1593 10999
rect 1593 10965 1627 10999
rect 1627 10965 1636 10999
rect 1584 10956 1636 10965
rect 8392 10999 8444 11008
rect 8392 10965 8401 10999
rect 8401 10965 8435 10999
rect 8435 10965 8444 10999
rect 8392 10956 8444 10965
rect 9312 11024 9364 11076
rect 10232 10956 10284 11008
rect 11060 11067 11112 11076
rect 11060 11033 11094 11067
rect 11094 11033 11112 11067
rect 13452 11092 13504 11144
rect 14280 11092 14332 11144
rect 14372 11135 14424 11144
rect 14372 11101 14381 11135
rect 14381 11101 14415 11135
rect 14415 11101 14424 11135
rect 14372 11092 14424 11101
rect 16120 11135 16172 11144
rect 16120 11101 16129 11135
rect 16129 11101 16163 11135
rect 16163 11101 16172 11135
rect 16120 11092 16172 11101
rect 16580 11092 16632 11144
rect 16764 11135 16816 11144
rect 16764 11101 16773 11135
rect 16773 11101 16807 11135
rect 16807 11101 16816 11135
rect 16764 11092 16816 11101
rect 20720 11169 20729 11203
rect 20729 11169 20763 11203
rect 20763 11169 20772 11203
rect 20720 11160 20772 11169
rect 18604 11092 18656 11144
rect 19432 11135 19484 11144
rect 19432 11101 19441 11135
rect 19441 11101 19475 11135
rect 19475 11101 19484 11135
rect 19432 11092 19484 11101
rect 20812 11092 20864 11144
rect 23480 11135 23532 11144
rect 23480 11101 23489 11135
rect 23489 11101 23523 11135
rect 23523 11101 23532 11135
rect 23480 11092 23532 11101
rect 23572 11092 23624 11144
rect 25688 11160 25740 11212
rect 24768 11135 24820 11144
rect 26240 11160 26292 11212
rect 26516 11160 26568 11212
rect 26608 11160 26660 11212
rect 24768 11101 24782 11135
rect 24782 11101 24816 11135
rect 24816 11101 24820 11135
rect 24768 11092 24820 11101
rect 11060 11024 11112 11033
rect 15476 11024 15528 11076
rect 16856 11024 16908 11076
rect 24584 11067 24636 11076
rect 24584 11033 24593 11067
rect 24593 11033 24627 11067
rect 24627 11033 24636 11067
rect 24584 11024 24636 11033
rect 25412 11024 25464 11076
rect 25964 11024 26016 11076
rect 26792 11135 26844 11144
rect 26792 11101 26801 11135
rect 26801 11101 26835 11135
rect 26835 11101 26844 11135
rect 26792 11092 26844 11101
rect 14096 10956 14148 11008
rect 15016 10956 15068 11008
rect 18236 10956 18288 11008
rect 21640 10956 21692 11008
rect 25596 10956 25648 11008
rect 26148 10956 26200 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 7564 10795 7616 10804
rect 7564 10761 7573 10795
rect 7573 10761 7607 10795
rect 7607 10761 7616 10795
rect 7564 10752 7616 10761
rect 9312 10684 9364 10736
rect 11060 10752 11112 10804
rect 15384 10795 15436 10804
rect 8208 10659 8260 10668
rect 8208 10625 8217 10659
rect 8217 10625 8251 10659
rect 8251 10625 8260 10659
rect 8208 10616 8260 10625
rect 9128 10616 9180 10668
rect 10784 10659 10836 10668
rect 10784 10625 10793 10659
rect 10793 10625 10827 10659
rect 10827 10625 10836 10659
rect 10784 10616 10836 10625
rect 11796 10659 11848 10668
rect 11796 10625 11805 10659
rect 11805 10625 11839 10659
rect 11839 10625 11848 10659
rect 11796 10616 11848 10625
rect 12256 10684 12308 10736
rect 12164 10659 12216 10668
rect 12164 10625 12173 10659
rect 12173 10625 12207 10659
rect 12207 10625 12216 10659
rect 15016 10684 15068 10736
rect 15384 10761 15393 10795
rect 15393 10761 15427 10795
rect 15427 10761 15436 10795
rect 15384 10752 15436 10761
rect 16120 10752 16172 10804
rect 16856 10795 16908 10804
rect 16856 10761 16865 10795
rect 16865 10761 16899 10795
rect 16899 10761 16908 10795
rect 16856 10752 16908 10761
rect 17960 10684 18012 10736
rect 19984 10752 20036 10804
rect 18420 10684 18472 10736
rect 12164 10616 12216 10625
rect 13176 10616 13228 10668
rect 14832 10616 14884 10668
rect 15476 10616 15528 10668
rect 15844 10659 15896 10668
rect 15844 10625 15853 10659
rect 15853 10625 15887 10659
rect 15887 10625 15896 10659
rect 15844 10616 15896 10625
rect 8484 10548 8536 10600
rect 10508 10548 10560 10600
rect 10692 10591 10744 10600
rect 10692 10557 10701 10591
rect 10701 10557 10735 10591
rect 10735 10557 10744 10591
rect 10692 10548 10744 10557
rect 14096 10548 14148 10600
rect 14740 10548 14792 10600
rect 18236 10659 18288 10668
rect 18236 10625 18271 10659
rect 18271 10625 18288 10659
rect 18236 10616 18288 10625
rect 20168 10616 20220 10668
rect 21272 10616 21324 10668
rect 21916 10616 21968 10668
rect 18144 10548 18196 10600
rect 18512 10548 18564 10600
rect 19892 10548 19944 10600
rect 21364 10548 21416 10600
rect 23572 10684 23624 10736
rect 22652 10591 22704 10600
rect 22652 10557 22661 10591
rect 22661 10557 22695 10591
rect 22695 10557 22704 10591
rect 22652 10548 22704 10557
rect 25688 10616 25740 10668
rect 26332 10659 26384 10668
rect 26332 10625 26341 10659
rect 26341 10625 26375 10659
rect 26375 10625 26384 10659
rect 26332 10616 26384 10625
rect 26516 10548 26568 10600
rect 9312 10412 9364 10464
rect 14188 10412 14240 10464
rect 14372 10412 14424 10464
rect 17960 10412 18012 10464
rect 24216 10480 24268 10532
rect 26148 10523 26200 10532
rect 26148 10489 26161 10523
rect 26161 10489 26195 10523
rect 26195 10489 26200 10523
rect 26148 10480 26200 10489
rect 20168 10412 20220 10464
rect 22284 10412 22336 10464
rect 22928 10412 22980 10464
rect 35808 10412 35860 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 8668 10208 8720 10260
rect 10508 10251 10560 10260
rect 8208 10140 8260 10192
rect 8024 10115 8076 10124
rect 8024 10081 8033 10115
rect 8033 10081 8067 10115
rect 8067 10081 8076 10115
rect 10508 10217 10517 10251
rect 10517 10217 10551 10251
rect 10551 10217 10560 10251
rect 10508 10208 10560 10217
rect 14832 10208 14884 10260
rect 16672 10208 16724 10260
rect 17960 10251 18012 10260
rect 15108 10140 15160 10192
rect 8024 10072 8076 10081
rect 8392 10004 8444 10056
rect 9312 10047 9364 10056
rect 9312 10013 9321 10047
rect 9321 10013 9355 10047
rect 9355 10013 9364 10047
rect 9312 10004 9364 10013
rect 9404 10004 9456 10056
rect 10324 10004 10376 10056
rect 10876 10004 10928 10056
rect 12256 10072 12308 10124
rect 11612 10004 11664 10056
rect 12900 10047 12952 10056
rect 12900 10013 12909 10047
rect 12909 10013 12943 10047
rect 12943 10013 12952 10047
rect 12900 10004 12952 10013
rect 14188 10047 14240 10056
rect 14188 10013 14197 10047
rect 14197 10013 14231 10047
rect 14231 10013 14240 10047
rect 14188 10004 14240 10013
rect 15200 10072 15252 10124
rect 14372 10004 14424 10056
rect 17960 10217 17969 10251
rect 17969 10217 18003 10251
rect 18003 10217 18012 10251
rect 17960 10208 18012 10217
rect 20168 10208 20220 10260
rect 22652 10208 22704 10260
rect 24584 10251 24636 10260
rect 24584 10217 24593 10251
rect 24593 10217 24627 10251
rect 24627 10217 24636 10251
rect 24584 10208 24636 10217
rect 25412 10251 25464 10260
rect 25412 10217 25421 10251
rect 25421 10217 25455 10251
rect 25455 10217 25464 10251
rect 25412 10208 25464 10217
rect 18052 10140 18104 10192
rect 24124 10140 24176 10192
rect 19064 10072 19116 10124
rect 20720 10072 20772 10124
rect 24676 10115 24728 10124
rect 24676 10081 24685 10115
rect 24685 10081 24719 10115
rect 24719 10081 24728 10115
rect 24676 10072 24728 10081
rect 17776 10047 17828 10056
rect 17776 10013 17785 10047
rect 17785 10013 17819 10047
rect 17819 10013 17828 10047
rect 17776 10004 17828 10013
rect 18604 10047 18656 10056
rect 18604 10013 18613 10047
rect 18613 10013 18647 10047
rect 18647 10013 18656 10047
rect 18604 10004 18656 10013
rect 19248 10047 19300 10056
rect 19248 10013 19257 10047
rect 19257 10013 19291 10047
rect 19291 10013 19300 10047
rect 19248 10004 19300 10013
rect 19340 10004 19392 10056
rect 25596 10072 25648 10124
rect 25320 10047 25372 10056
rect 25320 10013 25329 10047
rect 25329 10013 25363 10047
rect 25363 10013 25372 10047
rect 25320 10004 25372 10013
rect 25688 10004 25740 10056
rect 9128 9979 9180 9988
rect 9128 9945 9137 9979
rect 9137 9945 9171 9979
rect 9171 9945 9180 9979
rect 9128 9936 9180 9945
rect 10692 9936 10744 9988
rect 11336 9936 11388 9988
rect 15384 9936 15436 9988
rect 15936 9979 15988 9988
rect 15936 9945 15970 9979
rect 15970 9945 15988 9979
rect 15936 9936 15988 9945
rect 16580 9936 16632 9988
rect 22100 9936 22152 9988
rect 11520 9868 11572 9920
rect 12348 9911 12400 9920
rect 12348 9877 12357 9911
rect 12357 9877 12391 9911
rect 12391 9877 12400 9911
rect 12348 9868 12400 9877
rect 18420 9911 18472 9920
rect 18420 9877 18429 9911
rect 18429 9877 18463 9911
rect 18463 9877 18472 9911
rect 18420 9868 18472 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 9312 9664 9364 9716
rect 10692 9664 10744 9716
rect 11796 9664 11848 9716
rect 15936 9707 15988 9716
rect 15936 9673 15945 9707
rect 15945 9673 15979 9707
rect 15979 9673 15988 9707
rect 15936 9664 15988 9673
rect 10324 9596 10376 9648
rect 10876 9596 10928 9648
rect 9220 9571 9272 9580
rect 9220 9537 9229 9571
rect 9229 9537 9263 9571
rect 9263 9537 9272 9571
rect 9220 9528 9272 9537
rect 11336 9528 11388 9580
rect 11428 9528 11480 9580
rect 12256 9528 12308 9580
rect 13084 9528 13136 9580
rect 15384 9571 15436 9580
rect 11612 9503 11664 9512
rect 11612 9469 11621 9503
rect 11621 9469 11655 9503
rect 11655 9469 11664 9503
rect 11612 9460 11664 9469
rect 15384 9537 15393 9571
rect 15393 9537 15427 9571
rect 15427 9537 15436 9571
rect 15384 9528 15436 9537
rect 18420 9596 18472 9648
rect 19248 9596 19300 9648
rect 20720 9596 20772 9648
rect 15292 9460 15344 9512
rect 16212 9460 16264 9512
rect 20996 9528 21048 9580
rect 22744 9528 22796 9580
rect 16672 9503 16724 9512
rect 16672 9469 16681 9503
rect 16681 9469 16715 9503
rect 16715 9469 16724 9503
rect 16672 9460 16724 9469
rect 19064 9435 19116 9444
rect 19064 9401 19073 9435
rect 19073 9401 19107 9435
rect 19107 9401 19116 9435
rect 19064 9392 19116 9401
rect 11520 9367 11572 9376
rect 11520 9333 11529 9367
rect 11529 9333 11563 9367
rect 11563 9333 11572 9367
rect 11520 9324 11572 9333
rect 14740 9367 14792 9376
rect 14740 9333 14749 9367
rect 14749 9333 14783 9367
rect 14783 9333 14792 9367
rect 14740 9324 14792 9333
rect 21272 9367 21324 9376
rect 21272 9333 21281 9367
rect 21281 9333 21315 9367
rect 21315 9333 21324 9367
rect 21272 9324 21324 9333
rect 21364 9324 21416 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 9220 9120 9272 9172
rect 15016 9120 15068 9172
rect 18144 9120 18196 9172
rect 19432 9120 19484 9172
rect 20996 9163 21048 9172
rect 20996 9129 21005 9163
rect 21005 9129 21039 9163
rect 21039 9129 21048 9163
rect 20996 9120 21048 9129
rect 22100 9163 22152 9172
rect 22100 9129 22109 9163
rect 22109 9129 22143 9163
rect 22143 9129 22152 9163
rect 22100 9120 22152 9129
rect 22744 9163 22796 9172
rect 22744 9129 22753 9163
rect 22753 9129 22787 9163
rect 22787 9129 22796 9163
rect 22744 9120 22796 9129
rect 16672 9052 16724 9104
rect 17776 9052 17828 9104
rect 8024 9027 8076 9036
rect 8024 8993 8033 9027
rect 8033 8993 8067 9027
rect 8067 8993 8076 9027
rect 8024 8984 8076 8993
rect 12256 8984 12308 9036
rect 20168 9027 20220 9036
rect 20168 8993 20177 9027
rect 20177 8993 20211 9027
rect 20211 8993 20220 9027
rect 20168 8984 20220 8993
rect 8300 8916 8352 8968
rect 10324 8959 10376 8968
rect 10324 8925 10333 8959
rect 10333 8925 10367 8959
rect 10367 8925 10376 8959
rect 10324 8916 10376 8925
rect 12348 8959 12400 8968
rect 12348 8925 12357 8959
rect 12357 8925 12391 8959
rect 12391 8925 12400 8959
rect 12348 8916 12400 8925
rect 13544 8959 13596 8968
rect 13544 8925 13553 8959
rect 13553 8925 13587 8959
rect 13587 8925 13596 8959
rect 13544 8916 13596 8925
rect 13728 8916 13780 8968
rect 10232 8780 10284 8832
rect 10692 8848 10744 8900
rect 10876 8780 10928 8832
rect 12532 8823 12584 8832
rect 12532 8789 12541 8823
rect 12541 8789 12575 8823
rect 12575 8789 12584 8823
rect 12532 8780 12584 8789
rect 16212 8916 16264 8968
rect 19064 8916 19116 8968
rect 21916 8984 21968 9036
rect 22284 8959 22336 8968
rect 22284 8925 22293 8959
rect 22293 8925 22327 8959
rect 22327 8925 22336 8959
rect 22284 8916 22336 8925
rect 22928 8959 22980 8968
rect 22928 8925 22937 8959
rect 22937 8925 22971 8959
rect 22971 8925 22980 8959
rect 22928 8916 22980 8925
rect 18052 8848 18104 8900
rect 16764 8823 16816 8832
rect 16764 8789 16773 8823
rect 16773 8789 16807 8823
rect 16807 8789 16816 8823
rect 16764 8780 16816 8789
rect 21272 8848 21324 8900
rect 18604 8780 18656 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 8300 8576 8352 8628
rect 9128 8576 9180 8628
rect 10692 8619 10744 8628
rect 10692 8585 10701 8619
rect 10701 8585 10735 8619
rect 10735 8585 10744 8619
rect 10692 8576 10744 8585
rect 11520 8576 11572 8628
rect 13544 8576 13596 8628
rect 16672 8576 16724 8628
rect 10324 8508 10376 8560
rect 10232 8483 10284 8492
rect 10232 8449 10241 8483
rect 10241 8449 10275 8483
rect 10275 8449 10284 8483
rect 10232 8440 10284 8449
rect 11612 8440 11664 8492
rect 13728 8508 13780 8560
rect 11980 8483 12032 8492
rect 11980 8449 12014 8483
rect 12014 8449 12032 8483
rect 14740 8508 14792 8560
rect 16764 8508 16816 8560
rect 11980 8440 12032 8449
rect 15292 8440 15344 8492
rect 17592 8440 17644 8492
rect 10324 8372 10376 8424
rect 13728 8372 13780 8424
rect 16580 8304 16632 8356
rect 17316 8236 17368 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 11428 8032 11480 8084
rect 11612 8032 11664 8084
rect 11980 8032 12032 8084
rect 12256 8032 12308 8084
rect 17224 8032 17276 8084
rect 18604 8075 18656 8084
rect 18604 8041 18613 8075
rect 18613 8041 18647 8075
rect 18647 8041 18656 8075
rect 18604 8032 18656 8041
rect 11336 7939 11388 7948
rect 11336 7905 11345 7939
rect 11345 7905 11379 7939
rect 11379 7905 11388 7939
rect 11336 7896 11388 7905
rect 16580 7896 16632 7948
rect 10324 7828 10376 7880
rect 11520 7871 11572 7880
rect 11520 7837 11529 7871
rect 11529 7837 11563 7871
rect 11563 7837 11572 7871
rect 11520 7828 11572 7837
rect 12532 7828 12584 7880
rect 17316 7828 17368 7880
rect 9772 7803 9824 7812
rect 9772 7769 9806 7803
rect 9806 7769 9824 7803
rect 9772 7760 9824 7769
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 9772 7531 9824 7540
rect 9772 7497 9781 7531
rect 9781 7497 9815 7531
rect 9815 7497 9824 7531
rect 9772 7488 9824 7497
rect 17592 7531 17644 7540
rect 17592 7497 17601 7531
rect 17601 7497 17635 7531
rect 17635 7497 17644 7531
rect 17592 7488 17644 7497
rect 9956 7395 10008 7404
rect 9956 7361 9965 7395
rect 9965 7361 9999 7395
rect 9999 7361 10008 7395
rect 9956 7352 10008 7361
rect 17224 7395 17276 7404
rect 17224 7361 17233 7395
rect 17233 7361 17267 7395
rect 17267 7361 17276 7395
rect 17224 7352 17276 7361
rect 17408 7395 17460 7404
rect 17408 7361 17417 7395
rect 17417 7361 17451 7395
rect 17451 7361 17460 7395
rect 17408 7352 17460 7361
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 9220 6783 9272 6792
rect 9220 6749 9229 6783
rect 9229 6749 9263 6783
rect 9263 6749 9272 6783
rect 9220 6740 9272 6749
rect 9956 6808 10008 6860
rect 11336 6740 11388 6792
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 9220 2592 9272 2644
rect 11244 2592 11296 2644
rect 17408 2456 17460 2508
rect 20 2388 72 2440
rect 10324 2388 10376 2440
rect 26516 2388 26568 2440
rect 30932 2388 30984 2440
rect 37740 2388 37792 2440
rect 20628 2252 20680 2304
rect 38016 2295 38068 2304
rect 38016 2261 38025 2295
rect 38025 2261 38059 2295
rect 38059 2261 38068 2295
rect 38016 2252 38068 2261
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect 3238 39200 3294 40000
rect 13542 39200 13598 40000
rect 23846 39200 23902 40000
rect 34150 39200 34206 40000
rect 34256 39222 34468 39250
rect 3252 37126 3280 39200
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 3792 37256 3844 37262
rect 3792 37198 3844 37204
rect 3240 37120 3292 37126
rect 3240 37062 3292 37068
rect 1492 32904 1544 32910
rect 1492 32846 1544 32852
rect 1400 22024 1452 22030
rect 1400 21966 1452 21972
rect 1412 21865 1440 21966
rect 1398 21856 1454 21865
rect 1398 21791 1454 21800
rect 1504 12918 1532 32846
rect 1584 32768 1636 32774
rect 1582 32736 1584 32745
rect 1636 32736 1638 32745
rect 1582 32671 1638 32680
rect 3804 13734 3832 37198
rect 13556 37126 13584 39200
rect 23860 37262 23888 39200
rect 34164 39114 34192 39200
rect 34256 39114 34284 39222
rect 34164 39086 34284 39114
rect 25228 37460 25280 37466
rect 25228 37402 25280 37408
rect 24492 37392 24544 37398
rect 24492 37334 24544 37340
rect 14924 37256 14976 37262
rect 14924 37198 14976 37204
rect 23848 37256 23900 37262
rect 23848 37198 23900 37204
rect 13544 37120 13596 37126
rect 13544 37062 13596 37068
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 13820 28076 13872 28082
rect 13820 28018 13872 28024
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 13832 25770 13860 28018
rect 14280 28008 14332 28014
rect 14280 27950 14332 27956
rect 14292 27470 14320 27950
rect 14280 27464 14332 27470
rect 14280 27406 14332 27412
rect 14740 27464 14792 27470
rect 14740 27406 14792 27412
rect 14292 26926 14320 27406
rect 14648 26988 14700 26994
rect 14648 26930 14700 26936
rect 14280 26920 14332 26926
rect 14280 26862 14332 26868
rect 14292 26586 14320 26862
rect 14280 26580 14332 26586
rect 14280 26522 14332 26528
rect 14372 26376 14424 26382
rect 14372 26318 14424 26324
rect 14004 26308 14056 26314
rect 14004 26250 14056 26256
rect 13912 25900 13964 25906
rect 13912 25842 13964 25848
rect 13820 25764 13872 25770
rect 13820 25706 13872 25712
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 12992 24880 13044 24886
rect 12992 24822 13044 24828
rect 13820 24880 13872 24886
rect 13820 24822 13872 24828
rect 10048 24744 10100 24750
rect 10048 24686 10100 24692
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 8576 23792 8628 23798
rect 8576 23734 8628 23740
rect 8392 23724 8444 23730
rect 8392 23666 8444 23672
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 8404 23322 8432 23666
rect 8392 23316 8444 23322
rect 8392 23258 8444 23264
rect 8404 23118 8432 23258
rect 7012 23112 7064 23118
rect 7012 23054 7064 23060
rect 8392 23112 8444 23118
rect 8392 23054 8444 23060
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 7024 21486 7052 23054
rect 7932 21888 7984 21894
rect 7932 21830 7984 21836
rect 7012 21480 7064 21486
rect 7012 21422 7064 21428
rect 7288 21480 7340 21486
rect 7288 21422 7340 21428
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 7300 19446 7328 21422
rect 7748 20392 7800 20398
rect 7748 20334 7800 20340
rect 7760 20058 7788 20334
rect 7944 20058 7972 21830
rect 8588 21078 8616 23734
rect 9220 23724 9272 23730
rect 9220 23666 9272 23672
rect 9232 23322 9260 23666
rect 9312 23656 9364 23662
rect 9312 23598 9364 23604
rect 9220 23316 9272 23322
rect 9220 23258 9272 23264
rect 9036 23180 9088 23186
rect 9036 23122 9088 23128
rect 8944 23112 8996 23118
rect 8944 23054 8996 23060
rect 8956 22642 8984 23054
rect 9048 22642 9076 23122
rect 9324 22778 9352 23598
rect 9680 23520 9732 23526
rect 9680 23462 9732 23468
rect 9312 22772 9364 22778
rect 9312 22714 9364 22720
rect 8944 22636 8996 22642
rect 8944 22578 8996 22584
rect 9036 22636 9088 22642
rect 9036 22578 9088 22584
rect 8852 22568 8904 22574
rect 8852 22510 8904 22516
rect 8760 22432 8812 22438
rect 8760 22374 8812 22380
rect 8576 21072 8628 21078
rect 8576 21014 8628 21020
rect 8392 20800 8444 20806
rect 8392 20742 8444 20748
rect 8404 20466 8432 20742
rect 8392 20460 8444 20466
rect 8392 20402 8444 20408
rect 8300 20256 8352 20262
rect 8300 20198 8352 20204
rect 7748 20052 7800 20058
rect 7748 19994 7800 20000
rect 7932 20052 7984 20058
rect 7932 19994 7984 20000
rect 7944 19922 7972 19994
rect 7932 19916 7984 19922
rect 7932 19858 7984 19864
rect 7288 19440 7340 19446
rect 7288 19382 7340 19388
rect 8024 19372 8076 19378
rect 8024 19314 8076 19320
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 8036 18970 8064 19314
rect 8024 18964 8076 18970
rect 8024 18906 8076 18912
rect 8312 18766 8340 20198
rect 8404 19922 8432 20402
rect 8772 20398 8800 22374
rect 8864 22030 8892 22510
rect 9692 22438 9720 23462
rect 10060 22642 10088 24686
rect 10232 24268 10284 24274
rect 10232 24210 10284 24216
rect 10244 23662 10272 24210
rect 11612 24200 11664 24206
rect 11610 24168 11612 24177
rect 11888 24200 11940 24206
rect 11664 24168 11666 24177
rect 10324 24132 10376 24138
rect 11888 24142 11940 24148
rect 11610 24103 11666 24112
rect 10324 24074 10376 24080
rect 10336 23798 10364 24074
rect 10324 23792 10376 23798
rect 10324 23734 10376 23740
rect 10232 23656 10284 23662
rect 10232 23598 10284 23604
rect 10244 23526 10272 23598
rect 10232 23520 10284 23526
rect 10232 23462 10284 23468
rect 10232 23112 10284 23118
rect 10336 23100 10364 23734
rect 11152 23724 11204 23730
rect 11152 23666 11204 23672
rect 10508 23588 10560 23594
rect 10508 23530 10560 23536
rect 10284 23072 10364 23100
rect 10416 23112 10468 23118
rect 10232 23054 10284 23060
rect 10416 23054 10468 23060
rect 10428 22778 10456 23054
rect 10416 22772 10468 22778
rect 10416 22714 10468 22720
rect 10520 22642 10548 23530
rect 10600 23248 10652 23254
rect 10600 23190 10652 23196
rect 10612 23118 10640 23190
rect 11164 23186 11192 23666
rect 11152 23180 11204 23186
rect 11152 23122 11204 23128
rect 10600 23112 10652 23118
rect 10600 23054 10652 23060
rect 9864 22636 9916 22642
rect 9864 22578 9916 22584
rect 10048 22636 10100 22642
rect 10048 22578 10100 22584
rect 10508 22636 10560 22642
rect 10508 22578 10560 22584
rect 9680 22432 9732 22438
rect 9680 22374 9732 22380
rect 9692 22098 9720 22374
rect 9680 22092 9732 22098
rect 9680 22034 9732 22040
rect 8852 22024 8904 22030
rect 8852 21966 8904 21972
rect 8864 21690 8892 21966
rect 8852 21684 8904 21690
rect 8852 21626 8904 21632
rect 9692 21146 9720 22034
rect 9772 21616 9824 21622
rect 9772 21558 9824 21564
rect 9680 21140 9732 21146
rect 9680 21082 9732 21088
rect 9784 20942 9812 21558
rect 9876 21350 9904 22578
rect 9956 22092 10008 22098
rect 9956 22034 10008 22040
rect 9864 21344 9916 21350
rect 9864 21286 9916 21292
rect 9772 20936 9824 20942
rect 9772 20878 9824 20884
rect 9876 20874 9904 21286
rect 9968 21078 9996 22034
rect 10060 21690 10088 22578
rect 10048 21684 10100 21690
rect 10048 21626 10100 21632
rect 10232 21684 10284 21690
rect 10232 21626 10284 21632
rect 10140 21412 10192 21418
rect 10140 21354 10192 21360
rect 10152 21146 10180 21354
rect 10140 21140 10192 21146
rect 10140 21082 10192 21088
rect 9956 21072 10008 21078
rect 9956 21014 10008 21020
rect 10244 21010 10272 21626
rect 10612 21078 10640 23054
rect 11060 22976 11112 22982
rect 11060 22918 11112 22924
rect 11072 22642 11100 22918
rect 11060 22636 11112 22642
rect 11060 22578 11112 22584
rect 11164 22166 11192 23122
rect 11152 22160 11204 22166
rect 11152 22102 11204 22108
rect 10968 21956 11020 21962
rect 10968 21898 11020 21904
rect 10416 21072 10468 21078
rect 10416 21014 10468 21020
rect 10600 21072 10652 21078
rect 10600 21014 10652 21020
rect 10048 21004 10100 21010
rect 10048 20946 10100 20952
rect 10232 21004 10284 21010
rect 10232 20946 10284 20952
rect 9864 20868 9916 20874
rect 9864 20810 9916 20816
rect 9680 20800 9732 20806
rect 9680 20742 9732 20748
rect 9772 20800 9824 20806
rect 9772 20742 9824 20748
rect 9692 20466 9720 20742
rect 9680 20460 9732 20466
rect 9680 20402 9732 20408
rect 8760 20392 8812 20398
rect 8760 20334 8812 20340
rect 8392 19916 8444 19922
rect 8392 19858 8444 19864
rect 8772 19854 8800 20334
rect 9128 20256 9180 20262
rect 9128 20198 9180 20204
rect 9140 19990 9168 20198
rect 9128 19984 9180 19990
rect 9128 19926 9180 19932
rect 8760 19848 8812 19854
rect 8760 19790 8812 19796
rect 9140 19514 9168 19926
rect 9128 19508 9180 19514
rect 9128 19450 9180 19456
rect 9404 19440 9456 19446
rect 9404 19382 9456 19388
rect 9678 19408 9734 19417
rect 8300 18760 8352 18766
rect 8300 18702 8352 18708
rect 9416 18290 9444 19382
rect 9678 19343 9734 19352
rect 9692 18766 9720 19343
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 9784 18698 9812 20742
rect 10060 20534 10088 20946
rect 10324 20936 10376 20942
rect 10324 20878 10376 20884
rect 10048 20528 10100 20534
rect 10048 20470 10100 20476
rect 10060 19990 10088 20470
rect 10336 20466 10364 20878
rect 10428 20466 10456 21014
rect 10600 20936 10652 20942
rect 10600 20878 10652 20884
rect 10612 20602 10640 20878
rect 10980 20806 11008 21898
rect 11164 21486 11192 22102
rect 11624 22030 11652 24103
rect 11900 23866 11928 24142
rect 11888 23860 11940 23866
rect 11888 23802 11940 23808
rect 12716 23792 12768 23798
rect 12716 23734 12768 23740
rect 12072 23724 12124 23730
rect 12072 23666 12124 23672
rect 12532 23724 12584 23730
rect 12532 23666 12584 23672
rect 11980 23180 12032 23186
rect 11980 23122 12032 23128
rect 11992 22030 12020 23122
rect 12084 22778 12112 23666
rect 12348 23588 12400 23594
rect 12348 23530 12400 23536
rect 12256 23248 12308 23254
rect 12256 23190 12308 23196
rect 12072 22772 12124 22778
rect 12072 22714 12124 22720
rect 12072 22636 12124 22642
rect 12072 22578 12124 22584
rect 12084 22438 12112 22578
rect 12072 22432 12124 22438
rect 12072 22374 12124 22380
rect 11612 22024 11664 22030
rect 11612 21966 11664 21972
rect 11977 22024 12029 22030
rect 11977 21966 12029 21972
rect 11704 21888 11756 21894
rect 11704 21830 11756 21836
rect 11152 21480 11204 21486
rect 11152 21422 11204 21428
rect 11716 20942 11744 21830
rect 11796 21140 11848 21146
rect 11796 21082 11848 21088
rect 11336 20936 11388 20942
rect 11336 20878 11388 20884
rect 11704 20936 11756 20942
rect 11704 20878 11756 20884
rect 10968 20800 11020 20806
rect 10968 20742 11020 20748
rect 10600 20596 10652 20602
rect 10600 20538 10652 20544
rect 10324 20460 10376 20466
rect 10324 20402 10376 20408
rect 10416 20460 10468 20466
rect 10416 20402 10468 20408
rect 10968 20460 11020 20466
rect 10968 20402 11020 20408
rect 10048 19984 10100 19990
rect 10048 19926 10100 19932
rect 10336 19514 10364 20402
rect 10980 19990 11008 20402
rect 10968 19984 11020 19990
rect 10968 19926 11020 19932
rect 10416 19780 10468 19786
rect 10416 19722 10468 19728
rect 10428 19553 10456 19722
rect 10508 19712 10560 19718
rect 10508 19654 10560 19660
rect 10600 19712 10652 19718
rect 10600 19654 10652 19660
rect 10414 19544 10470 19553
rect 10324 19508 10376 19514
rect 10414 19479 10470 19488
rect 10324 19450 10376 19456
rect 10232 19440 10284 19446
rect 10232 19382 10284 19388
rect 10244 18834 10272 19382
rect 10324 19372 10376 19378
rect 10324 19314 10376 19320
rect 10336 18970 10364 19314
rect 10324 18964 10376 18970
rect 10324 18906 10376 18912
rect 10336 18850 10364 18906
rect 10232 18828 10284 18834
rect 10336 18822 10456 18850
rect 10232 18770 10284 18776
rect 10428 18766 10456 18822
rect 10416 18760 10468 18766
rect 10416 18702 10468 18708
rect 9772 18692 9824 18698
rect 9772 18634 9824 18640
rect 9404 18284 9456 18290
rect 9404 18226 9456 18232
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 9416 16658 9444 18226
rect 9784 17678 9812 18634
rect 10520 18358 10548 19654
rect 10612 19446 10640 19654
rect 10980 19446 11008 19926
rect 11348 19854 11376 20878
rect 11336 19848 11388 19854
rect 11336 19790 11388 19796
rect 11060 19712 11112 19718
rect 11060 19654 11112 19660
rect 10600 19440 10652 19446
rect 10598 19408 10600 19417
rect 10784 19440 10836 19446
rect 10652 19408 10654 19417
rect 10784 19382 10836 19388
rect 10968 19440 11020 19446
rect 10968 19382 11020 19388
rect 10598 19343 10654 19352
rect 10600 19304 10652 19310
rect 10600 19246 10652 19252
rect 10612 18970 10640 19246
rect 10796 19242 10824 19382
rect 10784 19236 10836 19242
rect 10784 19178 10836 19184
rect 10600 18964 10652 18970
rect 10600 18906 10652 18912
rect 10508 18352 10560 18358
rect 10508 18294 10560 18300
rect 10612 17882 10640 18906
rect 10784 18148 10836 18154
rect 10784 18090 10836 18096
rect 10600 17876 10652 17882
rect 10600 17818 10652 17824
rect 10796 17678 10824 18090
rect 11072 17882 11100 19654
rect 11244 18624 11296 18630
rect 11244 18566 11296 18572
rect 11060 17876 11112 17882
rect 11060 17818 11112 17824
rect 11256 17678 11284 18566
rect 9772 17672 9824 17678
rect 9772 17614 9824 17620
rect 10600 17672 10652 17678
rect 10600 17614 10652 17620
rect 10784 17672 10836 17678
rect 10784 17614 10836 17620
rect 11244 17672 11296 17678
rect 11244 17614 11296 17620
rect 10324 17196 10376 17202
rect 10324 17138 10376 17144
rect 9404 16652 9456 16658
rect 9404 16594 9456 16600
rect 9416 16182 9444 16594
rect 9588 16516 9640 16522
rect 9588 16458 9640 16464
rect 9404 16176 9456 16182
rect 9404 16118 9456 16124
rect 8300 16108 8352 16114
rect 8300 16050 8352 16056
rect 8576 16108 8628 16114
rect 8576 16050 8628 16056
rect 8852 16108 8904 16114
rect 8852 16050 8904 16056
rect 7748 15904 7800 15910
rect 7748 15846 7800 15852
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 7012 15564 7064 15570
rect 7012 15506 7064 15512
rect 6920 14816 6972 14822
rect 6920 14758 6972 14764
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 6932 14414 6960 14758
rect 7024 14618 7052 15506
rect 7760 15502 7788 15846
rect 7748 15496 7800 15502
rect 7748 15438 7800 15444
rect 8312 15162 8340 16050
rect 8588 15706 8616 16050
rect 8864 15706 8892 16050
rect 8576 15700 8628 15706
rect 8576 15642 8628 15648
rect 8852 15700 8904 15706
rect 8852 15642 8904 15648
rect 9128 15496 9180 15502
rect 9128 15438 9180 15444
rect 8392 15360 8444 15366
rect 8392 15302 8444 15308
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 8404 15094 8432 15302
rect 9140 15162 9168 15438
rect 9128 15156 9180 15162
rect 9128 15098 9180 15104
rect 8392 15088 8444 15094
rect 8392 15030 8444 15036
rect 9416 15026 9444 16118
rect 9600 15706 9628 16458
rect 9956 15904 10008 15910
rect 9956 15846 10008 15852
rect 9588 15700 9640 15706
rect 9588 15642 9640 15648
rect 9968 15570 9996 15846
rect 9956 15564 10008 15570
rect 9956 15506 10008 15512
rect 9772 15496 9824 15502
rect 9772 15438 9824 15444
rect 9864 15496 9916 15502
rect 9864 15438 9916 15444
rect 9588 15360 9640 15366
rect 9588 15302 9640 15308
rect 9404 15020 9456 15026
rect 9404 14962 9456 14968
rect 8024 14952 8076 14958
rect 8024 14894 8076 14900
rect 7012 14612 7064 14618
rect 7012 14554 7064 14560
rect 6920 14408 6972 14414
rect 6920 14350 6972 14356
rect 3792 13728 3844 13734
rect 3792 13670 3844 13676
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 7024 13394 7052 14554
rect 8036 13938 8064 14894
rect 9600 14618 9628 15302
rect 9784 14618 9812 15438
rect 9876 15026 9904 15438
rect 9968 15094 9996 15506
rect 10140 15428 10192 15434
rect 10140 15370 10192 15376
rect 9956 15088 10008 15094
rect 9956 15030 10008 15036
rect 9864 15020 9916 15026
rect 9864 14962 9916 14968
rect 9588 14612 9640 14618
rect 9588 14554 9640 14560
rect 9772 14612 9824 14618
rect 9772 14554 9824 14560
rect 9600 14346 9628 14554
rect 9968 14482 9996 15030
rect 9956 14476 10008 14482
rect 9956 14418 10008 14424
rect 9588 14340 9640 14346
rect 9588 14282 9640 14288
rect 8300 14272 8352 14278
rect 8300 14214 8352 14220
rect 9956 14272 10008 14278
rect 9956 14214 10008 14220
rect 8312 14006 8340 14214
rect 9968 14074 9996 14214
rect 9956 14068 10008 14074
rect 9956 14010 10008 14016
rect 8300 14000 8352 14006
rect 8300 13942 8352 13948
rect 9772 14000 9824 14006
rect 9772 13942 9824 13948
rect 8024 13932 8076 13938
rect 8024 13874 8076 13880
rect 8760 13932 8812 13938
rect 8760 13874 8812 13880
rect 9588 13932 9640 13938
rect 9588 13874 9640 13880
rect 9680 13932 9732 13938
rect 9680 13874 9732 13880
rect 8484 13864 8536 13870
rect 8484 13806 8536 13812
rect 7012 13388 7064 13394
rect 7012 13330 7064 13336
rect 1492 12912 1544 12918
rect 1492 12854 1544 12860
rect 7024 12850 7052 13330
rect 8496 13326 8524 13806
rect 8772 13530 8800 13874
rect 9128 13864 9180 13870
rect 9128 13806 9180 13812
rect 8760 13524 8812 13530
rect 8760 13466 8812 13472
rect 8484 13320 8536 13326
rect 8484 13262 8536 13268
rect 7012 12844 7064 12850
rect 7012 12786 7064 12792
rect 8116 12844 8168 12850
rect 8116 12786 8168 12792
rect 8852 12844 8904 12850
rect 8852 12786 8904 12792
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 8128 12306 8156 12786
rect 8864 12442 8892 12786
rect 8852 12436 8904 12442
rect 8852 12378 8904 12384
rect 8116 12300 8168 12306
rect 8116 12242 8168 12248
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 8128 11150 8156 12242
rect 9140 12238 9168 13806
rect 9600 13530 9628 13874
rect 9588 13524 9640 13530
rect 9588 13466 9640 13472
rect 9692 13394 9720 13874
rect 9680 13388 9732 13394
rect 9680 13330 9732 13336
rect 9692 12782 9720 13330
rect 9784 13258 9812 13942
rect 10152 13530 10180 15370
rect 10232 15020 10284 15026
rect 10232 14962 10284 14968
rect 10244 14074 10272 14962
rect 10232 14068 10284 14074
rect 10232 14010 10284 14016
rect 10232 13728 10284 13734
rect 10232 13670 10284 13676
rect 10244 13530 10272 13670
rect 10140 13524 10192 13530
rect 10140 13466 10192 13472
rect 10232 13524 10284 13530
rect 10232 13466 10284 13472
rect 9772 13252 9824 13258
rect 9772 13194 9824 13200
rect 9956 12844 10008 12850
rect 9956 12786 10008 12792
rect 9680 12776 9732 12782
rect 9680 12718 9732 12724
rect 9680 12640 9732 12646
rect 9680 12582 9732 12588
rect 9128 12232 9180 12238
rect 9128 12174 9180 12180
rect 9496 12164 9548 12170
rect 9496 12106 9548 12112
rect 9508 11898 9536 12106
rect 9496 11892 9548 11898
rect 9496 11834 9548 11840
rect 9692 11762 9720 12582
rect 9968 12481 9996 12786
rect 9954 12472 10010 12481
rect 9954 12407 10010 12416
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 9680 11756 9732 11762
rect 9680 11698 9732 11704
rect 8208 11688 8260 11694
rect 8208 11630 8260 11636
rect 8116 11144 8168 11150
rect 8116 11086 8168 11092
rect 7564 11076 7616 11082
rect 7564 11018 7616 11024
rect 1584 11008 1636 11014
rect 1582 10976 1584 10985
rect 1636 10976 1638 10985
rect 1582 10911 1638 10920
rect 7576 10810 7604 11018
rect 7564 10804 7616 10810
rect 7564 10746 7616 10752
rect 8220 10674 8248 11630
rect 8392 11008 8444 11014
rect 8392 10950 8444 10956
rect 8208 10668 8260 10674
rect 8208 10610 8260 10616
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 8220 10198 8248 10610
rect 8404 10554 8432 10950
rect 8484 10600 8536 10606
rect 8404 10548 8484 10554
rect 8404 10542 8536 10548
rect 8404 10526 8524 10542
rect 8208 10192 8260 10198
rect 8208 10134 8260 10140
rect 8024 10124 8076 10130
rect 8024 10066 8076 10072
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 8036 9042 8064 10066
rect 8404 10062 8432 10526
rect 8680 10266 8708 11698
rect 10336 11694 10364 17138
rect 10612 16794 10640 17614
rect 11348 17270 11376 19790
rect 11808 19334 11836 21082
rect 11992 20874 12020 21966
rect 11980 20868 12032 20874
rect 11980 20810 12032 20816
rect 11992 20330 12020 20810
rect 12084 20482 12112 22374
rect 12268 22030 12296 23190
rect 12360 22574 12388 23530
rect 12544 23338 12572 23666
rect 12452 23322 12572 23338
rect 12452 23316 12584 23322
rect 12452 23310 12532 23316
rect 12452 22642 12480 23310
rect 12532 23258 12584 23264
rect 12728 23118 12756 23734
rect 12808 23520 12860 23526
rect 12808 23462 12860 23468
rect 12716 23112 12768 23118
rect 12716 23054 12768 23060
rect 12624 22976 12676 22982
rect 12624 22918 12676 22924
rect 12440 22636 12492 22642
rect 12440 22578 12492 22584
rect 12348 22568 12400 22574
rect 12348 22510 12400 22516
rect 12256 22024 12308 22030
rect 12256 21966 12308 21972
rect 12360 21418 12388 22510
rect 12636 21690 12664 22918
rect 12728 22574 12756 23054
rect 12820 22642 12848 23462
rect 12900 23112 12952 23118
rect 12900 23054 12952 23060
rect 12912 22778 12940 23054
rect 12900 22772 12952 22778
rect 12900 22714 12952 22720
rect 12808 22636 12860 22642
rect 12808 22578 12860 22584
rect 12716 22568 12768 22574
rect 12716 22510 12768 22516
rect 12624 21684 12676 21690
rect 12624 21626 12676 21632
rect 12624 21548 12676 21554
rect 12624 21490 12676 21496
rect 12348 21412 12400 21418
rect 12348 21354 12400 21360
rect 12256 21344 12308 21350
rect 12256 21286 12308 21292
rect 12084 20454 12204 20482
rect 12176 20398 12204 20454
rect 12164 20392 12216 20398
rect 12164 20334 12216 20340
rect 11980 20324 12032 20330
rect 11980 20266 12032 20272
rect 11992 19922 12020 20266
rect 11980 19916 12032 19922
rect 11980 19858 12032 19864
rect 11992 19446 12020 19858
rect 11980 19440 12032 19446
rect 11980 19382 12032 19388
rect 11808 19306 11928 19334
rect 11900 18766 11928 19306
rect 11888 18760 11940 18766
rect 11888 18702 11940 18708
rect 11900 18290 11928 18702
rect 11888 18284 11940 18290
rect 11888 18226 11940 18232
rect 12176 17678 12204 20334
rect 12268 19310 12296 21286
rect 12360 19922 12388 21354
rect 12636 20806 12664 21490
rect 12808 21480 12860 21486
rect 12808 21422 12860 21428
rect 12820 21146 12848 21422
rect 12808 21140 12860 21146
rect 12808 21082 12860 21088
rect 12820 20874 12848 21082
rect 12808 20868 12860 20874
rect 12808 20810 12860 20816
rect 12624 20800 12676 20806
rect 12624 20742 12676 20748
rect 12636 19922 12664 20742
rect 12348 19916 12400 19922
rect 12348 19858 12400 19864
rect 12624 19916 12676 19922
rect 12624 19858 12676 19864
rect 12820 19854 12848 20810
rect 12808 19848 12860 19854
rect 12808 19790 12860 19796
rect 12624 19712 12676 19718
rect 12624 19654 12676 19660
rect 12346 19544 12402 19553
rect 12346 19479 12402 19488
rect 12360 19446 12388 19479
rect 12348 19440 12400 19446
rect 12348 19382 12400 19388
rect 12256 19304 12308 19310
rect 12256 19246 12308 19252
rect 12164 17672 12216 17678
rect 12164 17614 12216 17620
rect 12360 17338 12388 19382
rect 12440 19236 12492 19242
rect 12440 19178 12492 19184
rect 12452 18358 12480 19178
rect 12636 19174 12664 19654
rect 13004 19394 13032 24822
rect 13452 24064 13504 24070
rect 13452 24006 13504 24012
rect 13464 23730 13492 24006
rect 13452 23724 13504 23730
rect 13452 23666 13504 23672
rect 13636 23724 13688 23730
rect 13636 23666 13688 23672
rect 13084 23520 13136 23526
rect 13084 23462 13136 23468
rect 13096 22098 13124 23462
rect 13176 23112 13228 23118
rect 13176 23054 13228 23060
rect 13084 22092 13136 22098
rect 13084 22034 13136 22040
rect 13084 21888 13136 21894
rect 13084 21830 13136 21836
rect 13096 21146 13124 21830
rect 13188 21622 13216 23054
rect 13648 22574 13676 23666
rect 13636 22568 13688 22574
rect 13636 22510 13688 22516
rect 13360 21888 13412 21894
rect 13360 21830 13412 21836
rect 13176 21616 13228 21622
rect 13176 21558 13228 21564
rect 13084 21140 13136 21146
rect 13084 21082 13136 21088
rect 13188 21078 13216 21558
rect 13268 21548 13320 21554
rect 13268 21490 13320 21496
rect 13176 21072 13228 21078
rect 13176 21014 13228 21020
rect 13280 20602 13308 21490
rect 13372 21010 13400 21830
rect 13452 21684 13504 21690
rect 13452 21626 13504 21632
rect 13360 21004 13412 21010
rect 13360 20946 13412 20952
rect 13464 20874 13492 21626
rect 13452 20868 13504 20874
rect 13452 20810 13504 20816
rect 13268 20596 13320 20602
rect 13268 20538 13320 20544
rect 13464 19990 13492 20810
rect 13636 20800 13688 20806
rect 13636 20742 13688 20748
rect 13648 20398 13676 20742
rect 13636 20392 13688 20398
rect 13636 20334 13688 20340
rect 13452 19984 13504 19990
rect 13452 19926 13504 19932
rect 13832 19904 13860 24822
rect 13924 24342 13952 25842
rect 14016 25498 14044 26250
rect 14384 26042 14412 26318
rect 14660 26042 14688 26930
rect 14372 26036 14424 26042
rect 14372 25978 14424 25984
rect 14648 26036 14700 26042
rect 14648 25978 14700 25984
rect 14648 25900 14700 25906
rect 14648 25842 14700 25848
rect 14004 25492 14056 25498
rect 14004 25434 14056 25440
rect 14096 25288 14148 25294
rect 14096 25230 14148 25236
rect 14280 25288 14332 25294
rect 14280 25230 14332 25236
rect 13912 24336 13964 24342
rect 13912 24278 13964 24284
rect 14108 24274 14136 25230
rect 14292 24954 14320 25230
rect 14280 24948 14332 24954
rect 14280 24890 14332 24896
rect 14280 24812 14332 24818
rect 14280 24754 14332 24760
rect 14096 24268 14148 24274
rect 14096 24210 14148 24216
rect 14292 24138 14320 24754
rect 14660 24682 14688 25842
rect 14752 25498 14780 27406
rect 14740 25492 14792 25498
rect 14740 25434 14792 25440
rect 14648 24676 14700 24682
rect 14648 24618 14700 24624
rect 14280 24132 14332 24138
rect 14280 24074 14332 24080
rect 14292 23866 14320 24074
rect 14464 24064 14516 24070
rect 14464 24006 14516 24012
rect 14280 23860 14332 23866
rect 14280 23802 14332 23808
rect 14476 23730 14504 24006
rect 14556 23792 14608 23798
rect 14556 23734 14608 23740
rect 14464 23724 14516 23730
rect 14464 23666 14516 23672
rect 14280 22704 14332 22710
rect 14280 22646 14332 22652
rect 14096 22024 14148 22030
rect 14096 21966 14148 21972
rect 14108 20602 14136 21966
rect 14292 20806 14320 22646
rect 14372 22636 14424 22642
rect 14372 22578 14424 22584
rect 14384 21690 14412 22578
rect 14476 22234 14504 23666
rect 14568 22710 14596 23734
rect 14832 22976 14884 22982
rect 14832 22918 14884 22924
rect 14844 22710 14872 22918
rect 14556 22704 14608 22710
rect 14556 22646 14608 22652
rect 14832 22704 14884 22710
rect 14832 22646 14884 22652
rect 14464 22228 14516 22234
rect 14464 22170 14516 22176
rect 14372 21684 14424 21690
rect 14372 21626 14424 21632
rect 14384 21350 14412 21626
rect 14936 21486 14964 37198
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 24400 36848 24452 36854
rect 24400 36790 24452 36796
rect 24308 36780 24360 36786
rect 24308 36722 24360 36728
rect 24320 36106 24348 36722
rect 24412 36378 24440 36790
rect 24400 36372 24452 36378
rect 24400 36314 24452 36320
rect 24308 36100 24360 36106
rect 24308 36042 24360 36048
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 23756 35692 23808 35698
rect 23756 35634 23808 35640
rect 23664 35488 23716 35494
rect 23664 35430 23716 35436
rect 20168 35080 20220 35086
rect 20168 35022 20220 35028
rect 20444 35080 20496 35086
rect 20444 35022 20496 35028
rect 20812 35080 20864 35086
rect 20812 35022 20864 35028
rect 20996 35080 21048 35086
rect 20996 35022 21048 35028
rect 21824 35080 21876 35086
rect 21824 35022 21876 35028
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 19984 34604 20036 34610
rect 19984 34546 20036 34552
rect 19996 33998 20024 34546
rect 20076 34128 20128 34134
rect 20076 34070 20128 34076
rect 19248 33992 19300 33998
rect 19248 33934 19300 33940
rect 19984 33992 20036 33998
rect 19984 33934 20036 33940
rect 19260 33318 19288 33934
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 19432 33516 19484 33522
rect 19432 33458 19484 33464
rect 18328 33312 18380 33318
rect 18328 33254 18380 33260
rect 19248 33312 19300 33318
rect 19248 33254 19300 33260
rect 16764 32904 16816 32910
rect 16764 32846 16816 32852
rect 16856 32904 16908 32910
rect 16856 32846 16908 32852
rect 17224 32904 17276 32910
rect 17224 32846 17276 32852
rect 18052 32904 18104 32910
rect 18052 32846 18104 32852
rect 16776 32434 16804 32846
rect 16304 32428 16356 32434
rect 16304 32370 16356 32376
rect 16764 32428 16816 32434
rect 16764 32370 16816 32376
rect 15292 32360 15344 32366
rect 15292 32302 15344 32308
rect 15304 32026 15332 32302
rect 16316 32026 16344 32370
rect 15292 32020 15344 32026
rect 15292 31962 15344 31968
rect 16304 32020 16356 32026
rect 16304 31962 16356 31968
rect 15660 31884 15712 31890
rect 15660 31826 15712 31832
rect 16212 31884 16264 31890
rect 16212 31826 16264 31832
rect 15476 31816 15528 31822
rect 15476 31758 15528 31764
rect 15488 31482 15516 31758
rect 15476 31476 15528 31482
rect 15476 31418 15528 31424
rect 15292 31340 15344 31346
rect 15292 31282 15344 31288
rect 15200 31204 15252 31210
rect 15200 31146 15252 31152
rect 15212 30938 15240 31146
rect 15304 31142 15332 31282
rect 15292 31136 15344 31142
rect 15292 31078 15344 31084
rect 15200 30932 15252 30938
rect 15200 30874 15252 30880
rect 15672 30734 15700 31826
rect 16224 31754 16252 31826
rect 16776 31822 16804 32370
rect 16868 32298 16896 32846
rect 17236 32366 17264 32846
rect 17316 32768 17368 32774
rect 17316 32710 17368 32716
rect 17328 32434 17356 32710
rect 17316 32428 17368 32434
rect 17316 32370 17368 32376
rect 17224 32360 17276 32366
rect 17224 32302 17276 32308
rect 16856 32292 16908 32298
rect 16856 32234 16908 32240
rect 16868 31822 16896 32234
rect 17328 32026 17356 32370
rect 17316 32020 17368 32026
rect 17316 31962 17368 31968
rect 16764 31816 16816 31822
rect 16764 31758 16816 31764
rect 16856 31816 16908 31822
rect 16856 31758 16908 31764
rect 16028 31748 16080 31754
rect 16028 31690 16080 31696
rect 16132 31726 16252 31754
rect 15936 31680 15988 31686
rect 15936 31622 15988 31628
rect 15844 31272 15896 31278
rect 15844 31214 15896 31220
rect 15660 30728 15712 30734
rect 15660 30670 15712 30676
rect 15672 30326 15700 30670
rect 15856 30598 15884 31214
rect 15948 30734 15976 31622
rect 16040 31482 16068 31690
rect 16028 31476 16080 31482
rect 16028 31418 16080 31424
rect 16132 31362 16160 31726
rect 16040 31346 16160 31362
rect 16028 31340 16160 31346
rect 16080 31334 16160 31340
rect 16028 31282 16080 31288
rect 16040 30802 16068 31282
rect 16776 30938 16804 31758
rect 16868 31482 16896 31758
rect 17040 31748 17092 31754
rect 17040 31690 17092 31696
rect 16856 31476 16908 31482
rect 16856 31418 16908 31424
rect 17052 31346 17080 31690
rect 18064 31686 18092 32846
rect 18144 32768 18196 32774
rect 18144 32710 18196 32716
rect 18156 32434 18184 32710
rect 18144 32428 18196 32434
rect 18144 32370 18196 32376
rect 18052 31680 18104 31686
rect 18052 31622 18104 31628
rect 18236 31680 18288 31686
rect 18236 31622 18288 31628
rect 16856 31340 16908 31346
rect 16856 31282 16908 31288
rect 17040 31340 17092 31346
rect 17040 31282 17092 31288
rect 17868 31340 17920 31346
rect 17868 31282 17920 31288
rect 16764 30932 16816 30938
rect 16764 30874 16816 30880
rect 16868 30818 16896 31282
rect 16948 31136 17000 31142
rect 16948 31078 17000 31084
rect 16028 30796 16080 30802
rect 16028 30738 16080 30744
rect 16776 30790 16896 30818
rect 15936 30728 15988 30734
rect 15936 30670 15988 30676
rect 15844 30592 15896 30598
rect 15844 30534 15896 30540
rect 15660 30320 15712 30326
rect 15660 30262 15712 30268
rect 15856 30258 15884 30534
rect 15948 30394 15976 30670
rect 15936 30388 15988 30394
rect 15936 30330 15988 30336
rect 15844 30252 15896 30258
rect 15844 30194 15896 30200
rect 15856 29578 15884 30194
rect 16040 29714 16068 30738
rect 16580 30728 16632 30734
rect 16580 30670 16632 30676
rect 16592 30258 16620 30670
rect 16776 30666 16804 30790
rect 16764 30660 16816 30666
rect 16764 30602 16816 30608
rect 16580 30252 16632 30258
rect 16580 30194 16632 30200
rect 16776 30190 16804 30602
rect 16764 30184 16816 30190
rect 16764 30126 16816 30132
rect 16580 30048 16632 30054
rect 16580 29990 16632 29996
rect 16028 29708 16080 29714
rect 16028 29650 16080 29656
rect 16592 29646 16620 29990
rect 16580 29640 16632 29646
rect 16580 29582 16632 29588
rect 15476 29572 15528 29578
rect 15476 29514 15528 29520
rect 15844 29572 15896 29578
rect 15844 29514 15896 29520
rect 16120 29572 16172 29578
rect 16120 29514 16172 29520
rect 15488 28762 15516 29514
rect 15856 29238 15884 29514
rect 15844 29232 15896 29238
rect 15844 29174 15896 29180
rect 16132 29170 16160 29514
rect 16120 29164 16172 29170
rect 16120 29106 16172 29112
rect 16592 28762 16620 29582
rect 15476 28756 15528 28762
rect 15476 28698 15528 28704
rect 16580 28756 16632 28762
rect 16580 28698 16632 28704
rect 16028 28552 16080 28558
rect 16028 28494 16080 28500
rect 15936 27464 15988 27470
rect 15936 27406 15988 27412
rect 15948 27130 15976 27406
rect 15936 27124 15988 27130
rect 15936 27066 15988 27072
rect 15948 26994 15976 27066
rect 15936 26988 15988 26994
rect 15936 26930 15988 26936
rect 15292 26920 15344 26926
rect 15292 26862 15344 26868
rect 16040 26874 16068 28494
rect 16120 28484 16172 28490
rect 16120 28426 16172 28432
rect 16132 28218 16160 28426
rect 16120 28212 16172 28218
rect 16120 28154 16172 28160
rect 16776 27402 16804 30126
rect 16960 30122 16988 31078
rect 17592 30728 17644 30734
rect 17592 30670 17644 30676
rect 17040 30592 17092 30598
rect 17040 30534 17092 30540
rect 17052 30258 17080 30534
rect 17604 30258 17632 30670
rect 17776 30592 17828 30598
rect 17776 30534 17828 30540
rect 17040 30252 17092 30258
rect 17040 30194 17092 30200
rect 17592 30252 17644 30258
rect 17592 30194 17644 30200
rect 16948 30116 17000 30122
rect 16948 30058 17000 30064
rect 16960 29238 16988 30058
rect 17052 29850 17080 30194
rect 17040 29844 17092 29850
rect 17040 29786 17092 29792
rect 17408 29708 17460 29714
rect 17408 29650 17460 29656
rect 17420 29306 17448 29650
rect 17408 29300 17460 29306
rect 17408 29242 17460 29248
rect 16948 29232 17000 29238
rect 16948 29174 17000 29180
rect 17604 29170 17632 30194
rect 17788 30190 17816 30534
rect 17880 30394 17908 31282
rect 17960 31272 18012 31278
rect 17960 31214 18012 31220
rect 17972 30870 18000 31214
rect 18052 31204 18104 31210
rect 18052 31146 18104 31152
rect 17960 30864 18012 30870
rect 17960 30806 18012 30812
rect 18064 30734 18092 31146
rect 18144 31136 18196 31142
rect 18144 31078 18196 31084
rect 18156 30870 18184 31078
rect 18248 30938 18276 31622
rect 18340 31482 18368 33254
rect 19064 32564 19116 32570
rect 19064 32506 19116 32512
rect 18972 32428 19024 32434
rect 18972 32370 19024 32376
rect 18604 32224 18656 32230
rect 18604 32166 18656 32172
rect 18616 31890 18644 32166
rect 18788 31952 18840 31958
rect 18788 31894 18840 31900
rect 18604 31884 18656 31890
rect 18604 31826 18656 31832
rect 18800 31482 18828 31894
rect 18328 31476 18380 31482
rect 18328 31418 18380 31424
rect 18788 31476 18840 31482
rect 18788 31418 18840 31424
rect 18984 31346 19012 32370
rect 19076 31362 19104 32506
rect 19156 32428 19208 32434
rect 19156 32370 19208 32376
rect 19168 32314 19196 32370
rect 19168 32298 19288 32314
rect 19168 32292 19300 32298
rect 19168 32286 19248 32292
rect 19168 31754 19196 32286
rect 19248 32234 19300 32240
rect 19444 32230 19472 33458
rect 19996 33454 20024 33934
rect 20088 33522 20116 34070
rect 20180 33980 20208 35022
rect 20260 34944 20312 34950
rect 20260 34886 20312 34892
rect 20352 34944 20404 34950
rect 20352 34886 20404 34892
rect 20272 34610 20300 34886
rect 20260 34604 20312 34610
rect 20260 34546 20312 34552
rect 20364 34542 20392 34886
rect 20352 34536 20404 34542
rect 20352 34478 20404 34484
rect 20456 34354 20484 35022
rect 20824 34746 20852 35022
rect 20812 34740 20864 34746
rect 20812 34682 20864 34688
rect 20364 34326 20484 34354
rect 20260 33992 20312 33998
rect 20180 33952 20260 33980
rect 20260 33934 20312 33940
rect 20272 33522 20300 33934
rect 20364 33862 20392 34326
rect 21008 34066 21036 35022
rect 21836 34746 21864 35022
rect 21824 34740 21876 34746
rect 21824 34682 21876 34688
rect 23676 34610 23704 35430
rect 23768 35018 23796 35634
rect 24032 35624 24084 35630
rect 24032 35566 24084 35572
rect 23848 35556 23900 35562
rect 23848 35498 23900 35504
rect 23860 35086 23888 35498
rect 24044 35086 24072 35566
rect 23848 35080 23900 35086
rect 23848 35022 23900 35028
rect 24032 35080 24084 35086
rect 24032 35022 24084 35028
rect 23756 35012 23808 35018
rect 23756 34954 23808 34960
rect 21088 34604 21140 34610
rect 21088 34546 21140 34552
rect 23664 34604 23716 34610
rect 23664 34546 23716 34552
rect 21100 34202 21128 34546
rect 23768 34542 23796 34954
rect 23572 34536 23624 34542
rect 23572 34478 23624 34484
rect 23756 34536 23808 34542
rect 23756 34478 23808 34484
rect 22836 34468 22888 34474
rect 22836 34410 22888 34416
rect 21088 34196 21140 34202
rect 21088 34138 21140 34144
rect 20996 34060 21048 34066
rect 20996 34002 21048 34008
rect 20812 33992 20864 33998
rect 20812 33934 20864 33940
rect 20352 33856 20404 33862
rect 20352 33798 20404 33804
rect 20720 33856 20772 33862
rect 20720 33798 20772 33804
rect 20364 33522 20392 33798
rect 20076 33516 20128 33522
rect 20076 33458 20128 33464
rect 20260 33516 20312 33522
rect 20260 33458 20312 33464
rect 20352 33516 20404 33522
rect 20352 33458 20404 33464
rect 19984 33448 20036 33454
rect 19984 33390 20036 33396
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 19984 32360 20036 32366
rect 19984 32302 20036 32308
rect 19432 32224 19484 32230
rect 19432 32166 19484 32172
rect 19432 31816 19484 31822
rect 19352 31776 19432 31804
rect 19168 31726 19288 31754
rect 19260 31482 19288 31726
rect 19352 31482 19380 31776
rect 19432 31758 19484 31764
rect 19432 31680 19484 31686
rect 19432 31622 19484 31628
rect 19248 31476 19300 31482
rect 19248 31418 19300 31424
rect 19340 31476 19392 31482
rect 19340 31418 19392 31424
rect 19076 31346 19196 31362
rect 18512 31340 18564 31346
rect 18512 31282 18564 31288
rect 18972 31340 19024 31346
rect 19076 31340 19208 31346
rect 19076 31334 19156 31340
rect 18972 31282 19024 31288
rect 19156 31282 19208 31288
rect 18236 30932 18288 30938
rect 18236 30874 18288 30880
rect 18144 30864 18196 30870
rect 18144 30806 18196 30812
rect 18052 30728 18104 30734
rect 17972 30688 18052 30716
rect 17868 30388 17920 30394
rect 17868 30330 17920 30336
rect 17776 30184 17828 30190
rect 17776 30126 17828 30132
rect 17788 30054 17816 30126
rect 17776 30048 17828 30054
rect 17776 29990 17828 29996
rect 17788 29306 17816 29990
rect 17776 29300 17828 29306
rect 17776 29242 17828 29248
rect 17592 29164 17644 29170
rect 17592 29106 17644 29112
rect 17224 28756 17276 28762
rect 17224 28698 17276 28704
rect 16948 28552 17000 28558
rect 16948 28494 17000 28500
rect 16856 27872 16908 27878
rect 16856 27814 16908 27820
rect 16868 27402 16896 27814
rect 16960 27674 16988 28494
rect 17040 28144 17092 28150
rect 17040 28086 17092 28092
rect 17132 28144 17184 28150
rect 17132 28086 17184 28092
rect 16948 27668 17000 27674
rect 16948 27610 17000 27616
rect 16764 27396 16816 27402
rect 16764 27338 16816 27344
rect 16856 27396 16908 27402
rect 16856 27338 16908 27344
rect 16120 27328 16172 27334
rect 16120 27270 16172 27276
rect 16132 26994 16160 27270
rect 16120 26988 16172 26994
rect 16120 26930 16172 26936
rect 16764 26988 16816 26994
rect 16764 26930 16816 26936
rect 15304 26382 15332 26862
rect 16040 26846 16160 26874
rect 15476 26580 15528 26586
rect 15476 26522 15528 26528
rect 15488 26382 15516 26522
rect 15292 26376 15344 26382
rect 15292 26318 15344 26324
rect 15476 26376 15528 26382
rect 15476 26318 15528 26324
rect 15200 25968 15252 25974
rect 15200 25910 15252 25916
rect 15016 24880 15068 24886
rect 15016 24822 15068 24828
rect 15028 24750 15056 24822
rect 15212 24750 15240 25910
rect 15384 25900 15436 25906
rect 15384 25842 15436 25848
rect 15396 25498 15424 25842
rect 15488 25702 15516 26318
rect 16132 26314 16160 26846
rect 16672 26784 16724 26790
rect 16672 26726 16724 26732
rect 16684 26382 16712 26726
rect 16776 26586 16804 26930
rect 16868 26790 16896 27338
rect 17052 27334 17080 28086
rect 17144 27538 17172 28086
rect 17236 27878 17264 28698
rect 17224 27872 17276 27878
rect 17224 27814 17276 27820
rect 17132 27532 17184 27538
rect 17132 27474 17184 27480
rect 17236 27470 17264 27814
rect 17224 27464 17276 27470
rect 17224 27406 17276 27412
rect 17040 27328 17092 27334
rect 17040 27270 17092 27276
rect 17604 26790 17632 29106
rect 17788 27606 17816 29242
rect 17880 29170 17908 30330
rect 17972 29646 18000 30688
rect 18052 30670 18104 30676
rect 18052 30592 18104 30598
rect 18052 30534 18104 30540
rect 18064 29850 18092 30534
rect 18052 29844 18104 29850
rect 18052 29786 18104 29792
rect 18248 29646 18276 30874
rect 18328 30728 18380 30734
rect 18328 30670 18380 30676
rect 18340 30394 18368 30670
rect 18524 30546 18552 31282
rect 18604 30592 18656 30598
rect 18524 30540 18604 30546
rect 18524 30534 18656 30540
rect 18524 30518 18644 30534
rect 18524 30394 18552 30518
rect 18328 30388 18380 30394
rect 18328 30330 18380 30336
rect 18512 30388 18564 30394
rect 18512 30330 18564 30336
rect 19168 30190 19196 31282
rect 19260 30258 19288 31418
rect 19352 31260 19380 31418
rect 19444 31414 19472 31622
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 19432 31408 19484 31414
rect 19432 31350 19484 31356
rect 19352 31232 19472 31260
rect 19340 30660 19392 30666
rect 19340 30602 19392 30608
rect 19248 30252 19300 30258
rect 19248 30194 19300 30200
rect 19156 30184 19208 30190
rect 19156 30126 19208 30132
rect 17960 29640 18012 29646
rect 17960 29582 18012 29588
rect 18236 29640 18288 29646
rect 18236 29582 18288 29588
rect 17868 29164 17920 29170
rect 17868 29106 17920 29112
rect 18512 29164 18564 29170
rect 18512 29106 18564 29112
rect 18236 29096 18288 29102
rect 18236 29038 18288 29044
rect 18248 28218 18276 29038
rect 18420 28960 18472 28966
rect 18420 28902 18472 28908
rect 18432 28558 18460 28902
rect 18420 28552 18472 28558
rect 18420 28494 18472 28500
rect 18328 28484 18380 28490
rect 18328 28426 18380 28432
rect 18236 28212 18288 28218
rect 18236 28154 18288 28160
rect 18340 28082 18368 28426
rect 18328 28076 18380 28082
rect 18328 28018 18380 28024
rect 17776 27600 17828 27606
rect 17776 27542 17828 27548
rect 18052 27464 18104 27470
rect 18104 27412 18368 27418
rect 18052 27406 18368 27412
rect 18064 27390 18368 27406
rect 18052 27056 18104 27062
rect 18052 26998 18104 27004
rect 17960 26988 18012 26994
rect 17960 26930 18012 26936
rect 17972 26790 18000 26930
rect 16856 26784 16908 26790
rect 16856 26726 16908 26732
rect 17592 26784 17644 26790
rect 17592 26726 17644 26732
rect 17776 26784 17828 26790
rect 17776 26726 17828 26732
rect 17960 26784 18012 26790
rect 17960 26726 18012 26732
rect 17788 26586 17816 26726
rect 16764 26580 16816 26586
rect 16764 26522 16816 26528
rect 17776 26580 17828 26586
rect 17776 26522 17828 26528
rect 16672 26376 16724 26382
rect 16672 26318 16724 26324
rect 16120 26308 16172 26314
rect 16120 26250 16172 26256
rect 16132 26042 16160 26250
rect 17972 26042 18000 26726
rect 16120 26036 16172 26042
rect 16120 25978 16172 25984
rect 17960 26036 18012 26042
rect 17960 25978 18012 25984
rect 15752 25900 15804 25906
rect 15752 25842 15804 25848
rect 15476 25696 15528 25702
rect 15476 25638 15528 25644
rect 15384 25492 15436 25498
rect 15384 25434 15436 25440
rect 15488 25378 15516 25638
rect 15764 25498 15792 25842
rect 16396 25832 16448 25838
rect 16396 25774 16448 25780
rect 15752 25492 15804 25498
rect 15752 25434 15804 25440
rect 15396 25362 15516 25378
rect 16408 25362 16436 25774
rect 18064 25498 18092 26998
rect 18340 26858 18368 27390
rect 18524 27334 18552 29106
rect 18604 29096 18656 29102
rect 18604 29038 18656 29044
rect 18616 27538 18644 29038
rect 19168 28762 19196 30126
rect 19260 28966 19288 30194
rect 19352 29850 19380 30602
rect 19444 30258 19472 31232
rect 19996 31142 20024 32302
rect 20168 32224 20220 32230
rect 20168 32166 20220 32172
rect 20180 31754 20208 32166
rect 20168 31748 20220 31754
rect 20168 31690 20220 31696
rect 20076 31340 20128 31346
rect 20076 31282 20128 31288
rect 19984 31136 20036 31142
rect 19984 31078 20036 31084
rect 20088 30938 20116 31282
rect 20180 31278 20208 31690
rect 20272 31482 20300 33458
rect 20364 32026 20392 33458
rect 20444 33448 20496 33454
rect 20444 33390 20496 33396
rect 20352 32020 20404 32026
rect 20352 31962 20404 31968
rect 20456 31754 20484 33390
rect 20732 32910 20760 33798
rect 20824 33590 20852 33934
rect 21008 33658 21036 34002
rect 20996 33652 21048 33658
rect 20996 33594 21048 33600
rect 20812 33584 20864 33590
rect 20812 33526 20864 33532
rect 22192 33516 22244 33522
rect 22192 33458 22244 33464
rect 20812 33448 20864 33454
rect 20812 33390 20864 33396
rect 20824 33114 20852 33390
rect 21088 33312 21140 33318
rect 21088 33254 21140 33260
rect 20812 33108 20864 33114
rect 20812 33050 20864 33056
rect 20720 32904 20772 32910
rect 20720 32846 20772 32852
rect 20824 32502 20852 33050
rect 21100 32570 21128 33254
rect 22204 32910 22232 33458
rect 22848 33454 22876 34410
rect 23584 34066 23612 34478
rect 24032 34468 24084 34474
rect 24032 34410 24084 34416
rect 23572 34060 23624 34066
rect 23572 34002 23624 34008
rect 23480 33992 23532 33998
rect 23480 33934 23532 33940
rect 23756 33992 23808 33998
rect 23756 33934 23808 33940
rect 23492 33454 23520 33934
rect 22284 33448 22336 33454
rect 22284 33390 22336 33396
rect 22836 33448 22888 33454
rect 22836 33390 22888 33396
rect 23480 33448 23532 33454
rect 23480 33390 23532 33396
rect 22296 33046 22324 33390
rect 22284 33040 22336 33046
rect 22284 32982 22336 32988
rect 22192 32904 22244 32910
rect 22192 32846 22244 32852
rect 21916 32768 21968 32774
rect 21916 32710 21968 32716
rect 21088 32564 21140 32570
rect 21088 32506 21140 32512
rect 20812 32496 20864 32502
rect 20812 32438 20864 32444
rect 21100 31958 21128 32506
rect 21928 32230 21956 32710
rect 22284 32496 22336 32502
rect 22284 32438 22336 32444
rect 21916 32224 21968 32230
rect 21916 32166 21968 32172
rect 21088 31952 21140 31958
rect 21088 31894 21140 31900
rect 21928 31822 21956 32166
rect 22296 31890 22324 32438
rect 22848 32434 22876 33390
rect 23664 33312 23716 33318
rect 23664 33254 23716 33260
rect 23676 32910 23704 33254
rect 23768 33114 23796 33934
rect 23940 33924 23992 33930
rect 23940 33866 23992 33872
rect 23952 33522 23980 33866
rect 24044 33522 24072 34410
rect 24124 34060 24176 34066
rect 24124 34002 24176 34008
rect 24136 33590 24164 34002
rect 24124 33584 24176 33590
rect 24124 33526 24176 33532
rect 23940 33516 23992 33522
rect 23940 33458 23992 33464
rect 24032 33516 24084 33522
rect 24032 33458 24084 33464
rect 23756 33108 23808 33114
rect 23756 33050 23808 33056
rect 23756 32972 23808 32978
rect 23756 32914 23808 32920
rect 23664 32904 23716 32910
rect 23664 32846 23716 32852
rect 23204 32768 23256 32774
rect 23204 32710 23256 32716
rect 22836 32428 22888 32434
rect 22836 32370 22888 32376
rect 23020 32428 23072 32434
rect 23020 32370 23072 32376
rect 22284 31884 22336 31890
rect 22284 31826 22336 31832
rect 21088 31816 21140 31822
rect 21088 31758 21140 31764
rect 21916 31816 21968 31822
rect 21916 31758 21968 31764
rect 20456 31726 20668 31754
rect 20260 31476 20312 31482
rect 20260 31418 20312 31424
rect 20168 31272 20220 31278
rect 20168 31214 20220 31220
rect 20260 31204 20312 31210
rect 20260 31146 20312 31152
rect 20076 30932 20128 30938
rect 20076 30874 20128 30880
rect 19524 30728 19576 30734
rect 19522 30696 19524 30705
rect 19576 30696 19578 30705
rect 19522 30631 19578 30640
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 19432 30252 19484 30258
rect 19432 30194 19484 30200
rect 20272 30190 20300 31146
rect 20442 30696 20498 30705
rect 20442 30631 20498 30640
rect 20352 30252 20404 30258
rect 20352 30194 20404 30200
rect 20260 30184 20312 30190
rect 20260 30126 20312 30132
rect 19340 29844 19392 29850
rect 19340 29786 19392 29792
rect 20076 29844 20128 29850
rect 20076 29786 20128 29792
rect 19984 29504 20036 29510
rect 19984 29446 20036 29452
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 19996 29238 20024 29446
rect 19984 29232 20036 29238
rect 19984 29174 20036 29180
rect 20088 29170 20116 29786
rect 20260 29572 20312 29578
rect 20260 29514 20312 29520
rect 20168 29504 20220 29510
rect 20168 29446 20220 29452
rect 19708 29164 19760 29170
rect 19708 29106 19760 29112
rect 20076 29164 20128 29170
rect 20076 29106 20128 29112
rect 19248 28960 19300 28966
rect 19248 28902 19300 28908
rect 19156 28756 19208 28762
rect 19156 28698 19208 28704
rect 19340 28688 19392 28694
rect 19340 28630 19392 28636
rect 18972 28416 19024 28422
rect 18972 28358 19024 28364
rect 18984 28082 19012 28358
rect 19352 28150 19380 28630
rect 19720 28558 19748 29106
rect 20088 28994 20116 29106
rect 19904 28966 20116 28994
rect 19904 28762 19932 28966
rect 19892 28756 19944 28762
rect 19892 28698 19944 28704
rect 19984 28756 20036 28762
rect 19984 28698 20036 28704
rect 19800 28620 19852 28626
rect 19996 28608 20024 28698
rect 19852 28580 20024 28608
rect 19800 28562 19852 28568
rect 19432 28552 19484 28558
rect 19432 28494 19484 28500
rect 19708 28552 19760 28558
rect 20180 28506 20208 29446
rect 20272 29170 20300 29514
rect 20364 29170 20392 30194
rect 20260 29164 20312 29170
rect 20260 29106 20312 29112
rect 20352 29164 20404 29170
rect 20352 29106 20404 29112
rect 20272 28966 20300 29106
rect 20260 28960 20312 28966
rect 20260 28902 20312 28908
rect 20272 28694 20300 28902
rect 20260 28688 20312 28694
rect 20260 28630 20312 28636
rect 19708 28494 19760 28500
rect 19340 28144 19392 28150
rect 19340 28086 19392 28092
rect 18972 28076 19024 28082
rect 18972 28018 19024 28024
rect 19444 28014 19472 28494
rect 19812 28490 20208 28506
rect 19800 28484 20208 28490
rect 19852 28478 20208 28484
rect 19800 28426 19852 28432
rect 19984 28416 20036 28422
rect 19984 28358 20036 28364
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 19996 28082 20024 28358
rect 19984 28076 20036 28082
rect 19984 28018 20036 28024
rect 19432 28008 19484 28014
rect 19432 27950 19484 27956
rect 19708 28008 19760 28014
rect 19708 27950 19760 27956
rect 18696 27872 18748 27878
rect 18696 27814 18748 27820
rect 18604 27532 18656 27538
rect 18604 27474 18656 27480
rect 18512 27328 18564 27334
rect 18512 27270 18564 27276
rect 18144 26852 18196 26858
rect 18144 26794 18196 26800
rect 18328 26852 18380 26858
rect 18328 26794 18380 26800
rect 18156 25974 18184 26794
rect 18236 26784 18288 26790
rect 18236 26726 18288 26732
rect 18248 26450 18276 26726
rect 18236 26444 18288 26450
rect 18236 26386 18288 26392
rect 18144 25968 18196 25974
rect 18144 25910 18196 25916
rect 18052 25492 18104 25498
rect 18052 25434 18104 25440
rect 15384 25356 15516 25362
rect 15436 25350 15516 25356
rect 16396 25356 16448 25362
rect 15384 25298 15436 25304
rect 16396 25298 16448 25304
rect 15292 25288 15344 25294
rect 15292 25230 15344 25236
rect 15016 24744 15068 24750
rect 15016 24686 15068 24692
rect 15200 24744 15252 24750
rect 15200 24686 15252 24692
rect 15200 24608 15252 24614
rect 15200 24550 15252 24556
rect 15212 24342 15240 24550
rect 15304 24342 15332 25230
rect 15200 24336 15252 24342
rect 15200 24278 15252 24284
rect 15292 24336 15344 24342
rect 15292 24278 15344 24284
rect 15014 24168 15070 24177
rect 15014 24103 15016 24112
rect 15068 24103 15070 24112
rect 15016 24074 15068 24080
rect 15028 23322 15056 24074
rect 15108 24064 15160 24070
rect 15108 24006 15160 24012
rect 15120 23866 15148 24006
rect 15108 23860 15160 23866
rect 15108 23802 15160 23808
rect 15016 23316 15068 23322
rect 15016 23258 15068 23264
rect 15120 23254 15148 23802
rect 15212 23594 15240 24278
rect 15200 23588 15252 23594
rect 15200 23530 15252 23536
rect 15108 23248 15160 23254
rect 15108 23190 15160 23196
rect 15292 22500 15344 22506
rect 15292 22442 15344 22448
rect 15200 22160 15252 22166
rect 15200 22102 15252 22108
rect 15212 22030 15240 22102
rect 15200 22024 15252 22030
rect 15200 21966 15252 21972
rect 14924 21480 14976 21486
rect 14924 21422 14976 21428
rect 14372 21344 14424 21350
rect 14372 21286 14424 21292
rect 14372 20936 14424 20942
rect 14372 20878 14424 20884
rect 14280 20800 14332 20806
rect 14280 20742 14332 20748
rect 14096 20596 14148 20602
rect 14096 20538 14148 20544
rect 14292 20466 14320 20742
rect 14280 20460 14332 20466
rect 14280 20402 14332 20408
rect 14292 20346 14320 20402
rect 14200 20318 14320 20346
rect 13832 19876 13952 19904
rect 13452 19712 13504 19718
rect 13452 19654 13504 19660
rect 13004 19366 13400 19394
rect 13464 19378 13492 19654
rect 13924 19530 13952 19876
rect 13648 19502 13952 19530
rect 13648 19378 13676 19502
rect 13004 19360 13032 19366
rect 12912 19332 13032 19360
rect 12716 19304 12768 19310
rect 12912 19292 12940 19332
rect 12768 19264 12940 19292
rect 13176 19304 13228 19310
rect 12716 19246 12768 19252
rect 13176 19246 13228 19252
rect 12624 19168 12676 19174
rect 12624 19110 12676 19116
rect 12992 19168 13044 19174
rect 12992 19110 13044 19116
rect 12716 18692 12768 18698
rect 12716 18634 12768 18640
rect 12728 18426 12756 18634
rect 12716 18420 12768 18426
rect 12716 18362 12768 18368
rect 12440 18352 12492 18358
rect 12440 18294 12492 18300
rect 13004 18290 13032 19110
rect 13188 18290 13216 19246
rect 13372 19174 13400 19366
rect 13452 19372 13504 19378
rect 13452 19314 13504 19320
rect 13636 19372 13688 19378
rect 13636 19314 13688 19320
rect 13820 19372 13872 19378
rect 13820 19314 13872 19320
rect 13360 19168 13412 19174
rect 13360 19110 13412 19116
rect 13832 18970 13860 19314
rect 13924 18970 13952 19502
rect 13820 18964 13872 18970
rect 13820 18906 13872 18912
rect 13912 18964 13964 18970
rect 13912 18906 13964 18912
rect 13832 18358 13860 18906
rect 13924 18850 13952 18906
rect 13924 18822 14044 18850
rect 14016 18426 14044 18822
rect 14004 18420 14056 18426
rect 14004 18362 14056 18368
rect 13820 18352 13872 18358
rect 13820 18294 13872 18300
rect 12992 18284 13044 18290
rect 12992 18226 13044 18232
rect 13176 18284 13228 18290
rect 13176 18226 13228 18232
rect 12348 17332 12400 17338
rect 12348 17274 12400 17280
rect 14200 17270 14228 20318
rect 14384 19854 14412 20878
rect 15304 20602 15332 22442
rect 15396 22438 15424 25298
rect 16120 25288 16172 25294
rect 16120 25230 16172 25236
rect 16672 25288 16724 25294
rect 16672 25230 16724 25236
rect 17960 25288 18012 25294
rect 17960 25230 18012 25236
rect 15936 24812 15988 24818
rect 15936 24754 15988 24760
rect 15660 24132 15712 24138
rect 15660 24074 15712 24080
rect 15844 24132 15896 24138
rect 15844 24074 15896 24080
rect 15476 22636 15528 22642
rect 15476 22578 15528 22584
rect 15384 22432 15436 22438
rect 15384 22374 15436 22380
rect 15396 21962 15424 22374
rect 15488 22166 15516 22578
rect 15672 22574 15700 24074
rect 15660 22568 15712 22574
rect 15660 22510 15712 22516
rect 15672 22166 15700 22510
rect 15476 22160 15528 22166
rect 15476 22102 15528 22108
rect 15660 22160 15712 22166
rect 15660 22102 15712 22108
rect 15660 22024 15712 22030
rect 15856 22001 15884 24074
rect 15948 23866 15976 24754
rect 16132 24410 16160 25230
rect 16684 24682 16712 25230
rect 16764 24744 16816 24750
rect 16764 24686 16816 24692
rect 16672 24676 16724 24682
rect 16672 24618 16724 24624
rect 16120 24404 16172 24410
rect 16120 24346 16172 24352
rect 16488 24404 16540 24410
rect 16488 24346 16540 24352
rect 15936 23860 15988 23866
rect 15936 23802 15988 23808
rect 16396 23724 16448 23730
rect 16396 23666 16448 23672
rect 16408 22982 16436 23666
rect 16500 23526 16528 24346
rect 16776 24138 16804 24686
rect 17776 24608 17828 24614
rect 17776 24550 17828 24556
rect 17500 24200 17552 24206
rect 17500 24142 17552 24148
rect 16764 24132 16816 24138
rect 16764 24074 16816 24080
rect 16856 23656 16908 23662
rect 16856 23598 16908 23604
rect 16488 23520 16540 23526
rect 16488 23462 16540 23468
rect 16396 22976 16448 22982
rect 16396 22918 16448 22924
rect 16408 22642 16436 22918
rect 16396 22636 16448 22642
rect 16396 22578 16448 22584
rect 16408 22098 16436 22578
rect 16500 22438 16528 23462
rect 16764 23112 16816 23118
rect 16764 23054 16816 23060
rect 16776 22778 16804 23054
rect 16764 22772 16816 22778
rect 16764 22714 16816 22720
rect 16488 22432 16540 22438
rect 16488 22374 16540 22380
rect 16396 22092 16448 22098
rect 16396 22034 16448 22040
rect 15936 22024 15988 22030
rect 15660 21966 15712 21972
rect 15842 21992 15898 22001
rect 15384 21956 15436 21962
rect 15384 21898 15436 21904
rect 15384 21616 15436 21622
rect 15382 21584 15384 21593
rect 15436 21584 15438 21593
rect 15382 21519 15438 21528
rect 15476 21548 15528 21554
rect 15476 21490 15528 21496
rect 15488 21350 15516 21490
rect 15476 21344 15528 21350
rect 15476 21286 15528 21292
rect 15672 21078 15700 21966
rect 15936 21966 15988 21972
rect 15842 21927 15898 21936
rect 15660 21072 15712 21078
rect 15660 21014 15712 21020
rect 15292 20596 15344 20602
rect 15292 20538 15344 20544
rect 15660 20392 15712 20398
rect 15660 20334 15712 20340
rect 14372 19848 14424 19854
rect 14372 19790 14424 19796
rect 14280 19780 14332 19786
rect 14280 19722 14332 19728
rect 14292 17882 14320 19722
rect 14384 18766 14412 19790
rect 15672 19718 15700 20334
rect 15856 20262 15884 21927
rect 15948 21554 15976 21966
rect 16304 21888 16356 21894
rect 16304 21830 16356 21836
rect 15936 21548 15988 21554
rect 15936 21490 15988 21496
rect 16120 21548 16172 21554
rect 16120 21490 16172 21496
rect 15948 20806 15976 21490
rect 15936 20800 15988 20806
rect 15936 20742 15988 20748
rect 15844 20256 15896 20262
rect 15844 20198 15896 20204
rect 16132 19922 16160 21490
rect 16212 21072 16264 21078
rect 16212 21014 16264 21020
rect 16120 19916 16172 19922
rect 16120 19858 16172 19864
rect 15844 19848 15896 19854
rect 15844 19790 15896 19796
rect 15660 19712 15712 19718
rect 15660 19654 15712 19660
rect 15384 19372 15436 19378
rect 15384 19314 15436 19320
rect 15016 19168 15068 19174
rect 15016 19110 15068 19116
rect 15108 19168 15160 19174
rect 15108 19110 15160 19116
rect 14372 18760 14424 18766
rect 14372 18702 14424 18708
rect 14280 17876 14332 17882
rect 14280 17818 14332 17824
rect 15028 17678 15056 19110
rect 15120 18970 15148 19110
rect 15396 18970 15424 19314
rect 15672 19310 15700 19654
rect 15660 19304 15712 19310
rect 15660 19246 15712 19252
rect 15108 18964 15160 18970
rect 15108 18906 15160 18912
rect 15384 18964 15436 18970
rect 15384 18906 15436 18912
rect 15290 18728 15346 18737
rect 15290 18663 15346 18672
rect 15304 18290 15332 18663
rect 15292 18284 15344 18290
rect 15292 18226 15344 18232
rect 15856 17746 15884 19790
rect 15936 19508 15988 19514
rect 15936 19450 15988 19456
rect 15948 18358 15976 19450
rect 15936 18352 15988 18358
rect 15936 18294 15988 18300
rect 16224 17746 16252 21014
rect 16316 18698 16344 21830
rect 16868 21468 16896 23598
rect 17040 22568 17092 22574
rect 17040 22510 17092 22516
rect 17052 21978 17080 22510
rect 16960 21962 17080 21978
rect 16948 21956 17080 21962
rect 17000 21950 17080 21956
rect 16948 21898 17000 21904
rect 16776 21440 16896 21468
rect 16580 21344 16632 21350
rect 16580 21286 16632 21292
rect 16488 21140 16540 21146
rect 16488 21082 16540 21088
rect 16396 20392 16448 20398
rect 16396 20334 16448 20340
rect 16408 19334 16436 20334
rect 16500 19922 16528 21082
rect 16592 20330 16620 21286
rect 16580 20324 16632 20330
rect 16580 20266 16632 20272
rect 16488 19916 16540 19922
rect 16488 19858 16540 19864
rect 16500 19514 16528 19858
rect 16488 19508 16540 19514
rect 16488 19450 16540 19456
rect 16408 19306 16528 19334
rect 16396 18760 16448 18766
rect 16396 18702 16448 18708
rect 16304 18692 16356 18698
rect 16304 18634 16356 18640
rect 16408 18222 16436 18702
rect 16500 18290 16528 19306
rect 16776 19242 16804 21440
rect 16960 21146 16988 21898
rect 17132 21888 17184 21894
rect 17052 21836 17132 21842
rect 17052 21830 17184 21836
rect 17052 21814 17172 21830
rect 16948 21140 17000 21146
rect 16948 21082 17000 21088
rect 16856 20256 16908 20262
rect 16856 20198 16908 20204
rect 16764 19236 16816 19242
rect 16764 19178 16816 19184
rect 16776 18970 16804 19178
rect 16764 18964 16816 18970
rect 16764 18906 16816 18912
rect 16580 18692 16632 18698
rect 16580 18634 16632 18640
rect 16764 18692 16816 18698
rect 16764 18634 16816 18640
rect 16592 18426 16620 18634
rect 16580 18420 16632 18426
rect 16580 18362 16632 18368
rect 16488 18284 16540 18290
rect 16488 18226 16540 18232
rect 16396 18216 16448 18222
rect 16396 18158 16448 18164
rect 15844 17740 15896 17746
rect 15844 17682 15896 17688
rect 16212 17740 16264 17746
rect 16212 17682 16264 17688
rect 15016 17672 15068 17678
rect 15016 17614 15068 17620
rect 14924 17536 14976 17542
rect 14924 17478 14976 17484
rect 11336 17264 11388 17270
rect 11336 17206 11388 17212
rect 12808 17264 12860 17270
rect 12808 17206 12860 17212
rect 14188 17264 14240 17270
rect 14188 17206 14240 17212
rect 12716 17196 12768 17202
rect 12716 17138 12768 17144
rect 12624 16992 12676 16998
rect 12624 16934 12676 16940
rect 10600 16788 10652 16794
rect 10600 16730 10652 16736
rect 12636 16590 12664 16934
rect 12728 16726 12756 17138
rect 12820 16794 12848 17206
rect 12900 17196 12952 17202
rect 12900 17138 12952 17144
rect 14096 17196 14148 17202
rect 14096 17138 14148 17144
rect 14740 17196 14792 17202
rect 14740 17138 14792 17144
rect 12808 16788 12860 16794
rect 12808 16730 12860 16736
rect 12716 16720 12768 16726
rect 12716 16662 12768 16668
rect 12912 16590 12940 17138
rect 13084 17128 13136 17134
rect 13084 17070 13136 17076
rect 13096 16658 13124 17070
rect 13084 16652 13136 16658
rect 13084 16594 13136 16600
rect 12624 16584 12676 16590
rect 12624 16526 12676 16532
rect 12900 16584 12952 16590
rect 12900 16526 12952 16532
rect 11796 16448 11848 16454
rect 11796 16390 11848 16396
rect 11808 15978 11836 16390
rect 12636 16250 12664 16526
rect 12624 16244 12676 16250
rect 12624 16186 12676 16192
rect 12256 16040 12308 16046
rect 12256 15982 12308 15988
rect 11796 15972 11848 15978
rect 11796 15914 11848 15920
rect 11808 15570 11836 15914
rect 12268 15638 12296 15982
rect 12912 15706 12940 16526
rect 12900 15700 12952 15706
rect 12900 15642 12952 15648
rect 12256 15632 12308 15638
rect 12256 15574 12308 15580
rect 11796 15564 11848 15570
rect 11796 15506 11848 15512
rect 10876 15496 10928 15502
rect 10876 15438 10928 15444
rect 11336 15496 11388 15502
rect 11336 15438 11388 15444
rect 10600 14952 10652 14958
rect 10600 14894 10652 14900
rect 10612 14618 10640 14894
rect 10888 14618 10916 15438
rect 10968 14816 11020 14822
rect 10968 14758 11020 14764
rect 10600 14612 10652 14618
rect 10600 14554 10652 14560
rect 10876 14612 10928 14618
rect 10876 14554 10928 14560
rect 10980 14414 11008 14758
rect 11060 14476 11112 14482
rect 11060 14418 11112 14424
rect 10968 14408 11020 14414
rect 10968 14350 11020 14356
rect 10968 13252 11020 13258
rect 10968 13194 11020 13200
rect 10980 12442 11008 13194
rect 11072 12714 11100 14418
rect 11060 12708 11112 12714
rect 11060 12650 11112 12656
rect 10968 12436 11020 12442
rect 10968 12378 11020 12384
rect 11244 12164 11296 12170
rect 11244 12106 11296 12112
rect 10324 11688 10376 11694
rect 10324 11630 10376 11636
rect 9036 11552 9088 11558
rect 9036 11494 9088 11500
rect 9048 11150 9076 11494
rect 9036 11144 9088 11150
rect 9036 11086 9088 11092
rect 10232 11144 10284 11150
rect 10232 11086 10284 11092
rect 10876 11144 10928 11150
rect 10876 11086 10928 11092
rect 9312 11076 9364 11082
rect 9312 11018 9364 11024
rect 9324 10742 9352 11018
rect 10244 11014 10272 11086
rect 10232 11008 10284 11014
rect 10232 10950 10284 10956
rect 9312 10736 9364 10742
rect 9312 10678 9364 10684
rect 9128 10668 9180 10674
rect 9128 10610 9180 10616
rect 8668 10260 8720 10266
rect 8668 10202 8720 10208
rect 8392 10056 8444 10062
rect 8392 9998 8444 10004
rect 9140 9994 9168 10610
rect 9324 10554 9352 10678
rect 10784 10668 10836 10674
rect 10784 10610 10836 10616
rect 10508 10600 10560 10606
rect 9324 10526 9444 10554
rect 10508 10542 10560 10548
rect 10692 10600 10744 10606
rect 10692 10542 10744 10548
rect 9312 10464 9364 10470
rect 9312 10406 9364 10412
rect 9324 10062 9352 10406
rect 9416 10062 9444 10526
rect 10520 10266 10548 10542
rect 10508 10260 10560 10266
rect 10508 10202 10560 10208
rect 9312 10056 9364 10062
rect 9312 9998 9364 10004
rect 9404 10056 9456 10062
rect 9404 9998 9456 10004
rect 10324 10056 10376 10062
rect 10324 9998 10376 10004
rect 9128 9988 9180 9994
rect 9128 9930 9180 9936
rect 8024 9036 8076 9042
rect 8024 8978 8076 8984
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 8312 8634 8340 8910
rect 9140 8634 9168 9930
rect 9324 9722 9352 9998
rect 9312 9716 9364 9722
rect 9312 9658 9364 9664
rect 10336 9654 10364 9998
rect 10704 9994 10732 10542
rect 10692 9988 10744 9994
rect 10692 9930 10744 9936
rect 10704 9722 10732 9930
rect 10796 9738 10824 10610
rect 10888 10062 10916 11086
rect 11060 11076 11112 11082
rect 11060 11018 11112 11024
rect 11072 10810 11100 11018
rect 11060 10804 11112 10810
rect 11060 10746 11112 10752
rect 10876 10056 10928 10062
rect 10876 9998 10928 10004
rect 10692 9716 10744 9722
rect 10796 9710 10916 9738
rect 10692 9658 10744 9664
rect 10888 9654 10916 9710
rect 10324 9648 10376 9654
rect 10324 9590 10376 9596
rect 10876 9648 10928 9654
rect 10876 9590 10928 9596
rect 9220 9580 9272 9586
rect 9220 9522 9272 9528
rect 9232 9178 9260 9522
rect 9220 9172 9272 9178
rect 9220 9114 9272 9120
rect 10336 8974 10364 9590
rect 10324 8968 10376 8974
rect 10324 8910 10376 8916
rect 10232 8832 10284 8838
rect 10232 8774 10284 8780
rect 8300 8628 8352 8634
rect 8300 8570 8352 8576
rect 9128 8628 9180 8634
rect 9128 8570 9180 8576
rect 10244 8498 10272 8774
rect 10336 8566 10364 8910
rect 10692 8900 10744 8906
rect 10692 8842 10744 8848
rect 10704 8634 10732 8842
rect 10888 8838 10916 9590
rect 10876 8832 10928 8838
rect 10876 8774 10928 8780
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 10324 8560 10376 8566
rect 10324 8502 10376 8508
rect 10232 8492 10284 8498
rect 10232 8434 10284 8440
rect 10336 8430 10364 8502
rect 10324 8424 10376 8430
rect 10324 8366 10376 8372
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 10336 7886 10364 8366
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 9772 7812 9824 7818
rect 9772 7754 9824 7760
rect 9784 7546 9812 7754
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 9956 7404 10008 7410
rect 9956 7346 10008 7352
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 9968 6866 9996 7346
rect 9956 6860 10008 6866
rect 9956 6802 10008 6808
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 9232 2650 9260 6734
rect 11256 2650 11284 12106
rect 11348 11558 11376 15438
rect 11704 14816 11756 14822
rect 11704 14758 11756 14764
rect 11520 14340 11572 14346
rect 11520 14282 11572 14288
rect 11532 12782 11560 14282
rect 11612 14000 11664 14006
rect 11612 13942 11664 13948
rect 11624 13326 11652 13942
rect 11716 13938 11744 14758
rect 11704 13932 11756 13938
rect 11704 13874 11756 13880
rect 11796 13796 11848 13802
rect 11796 13738 11848 13744
rect 11612 13320 11664 13326
rect 11612 13262 11664 13268
rect 11808 13258 11836 13738
rect 11796 13252 11848 13258
rect 11796 13194 11848 13200
rect 11612 12844 11664 12850
rect 11612 12786 11664 12792
rect 11520 12776 11572 12782
rect 11520 12718 11572 12724
rect 11624 12374 11652 12786
rect 11612 12368 11664 12374
rect 11612 12310 11664 12316
rect 11808 12306 11836 13194
rect 12268 12306 12296 15574
rect 12440 15088 12492 15094
rect 12440 15030 12492 15036
rect 12452 14414 12480 15030
rect 12716 15020 12768 15026
rect 12716 14962 12768 14968
rect 12440 14408 12492 14414
rect 12440 14350 12492 14356
rect 12728 14074 12756 14962
rect 13096 14618 13124 16594
rect 14108 16590 14136 17138
rect 14188 17128 14240 17134
rect 14188 17070 14240 17076
rect 14200 16794 14228 17070
rect 14188 16788 14240 16794
rect 14188 16730 14240 16736
rect 13544 16584 13596 16590
rect 13544 16526 13596 16532
rect 14096 16584 14148 16590
rect 14096 16526 14148 16532
rect 13360 16448 13412 16454
rect 13360 16390 13412 16396
rect 13372 16182 13400 16390
rect 13360 16176 13412 16182
rect 13360 16118 13412 16124
rect 13176 16108 13228 16114
rect 13176 16050 13228 16056
rect 13188 14958 13216 16050
rect 13556 15706 13584 16526
rect 14108 16250 14136 16526
rect 14096 16244 14148 16250
rect 14096 16186 14148 16192
rect 14200 16114 14228 16730
rect 14752 16726 14780 17138
rect 14740 16720 14792 16726
rect 14740 16662 14792 16668
rect 14936 16590 14964 17478
rect 14924 16584 14976 16590
rect 14924 16526 14976 16532
rect 14188 16108 14240 16114
rect 14188 16050 14240 16056
rect 13544 15700 13596 15706
rect 13544 15642 13596 15648
rect 13452 15496 13504 15502
rect 13452 15438 13504 15444
rect 15016 15496 15068 15502
rect 15016 15438 15068 15444
rect 13176 14952 13228 14958
rect 13176 14894 13228 14900
rect 13084 14612 13136 14618
rect 13084 14554 13136 14560
rect 12900 14408 12952 14414
rect 12900 14350 12952 14356
rect 12716 14068 12768 14074
rect 12716 14010 12768 14016
rect 12912 13938 12940 14350
rect 13188 14346 13216 14894
rect 13176 14340 13228 14346
rect 13176 14282 13228 14288
rect 12624 13932 12676 13938
rect 12624 13874 12676 13880
rect 12900 13932 12952 13938
rect 12900 13874 12952 13880
rect 12532 13184 12584 13190
rect 12532 13126 12584 13132
rect 12544 12918 12572 13126
rect 12532 12912 12584 12918
rect 12532 12854 12584 12860
rect 12348 12844 12400 12850
rect 12348 12786 12400 12792
rect 12360 12730 12388 12786
rect 12360 12702 12480 12730
rect 12452 12442 12480 12702
rect 12440 12436 12492 12442
rect 12440 12378 12492 12384
rect 11796 12300 11848 12306
rect 11796 12242 11848 12248
rect 12256 12300 12308 12306
rect 12256 12242 12308 12248
rect 11336 11552 11388 11558
rect 11336 11494 11388 11500
rect 12164 11552 12216 11558
rect 12164 11494 12216 11500
rect 12176 10674 12204 11494
rect 12268 11354 12296 12242
rect 12636 11762 12664 13874
rect 13188 12782 13216 14282
rect 13464 13938 13492 15438
rect 14556 14816 14608 14822
rect 14556 14758 14608 14764
rect 14568 14482 14596 14758
rect 14556 14476 14608 14482
rect 14556 14418 14608 14424
rect 15028 14414 15056 15438
rect 15200 15360 15252 15366
rect 15200 15302 15252 15308
rect 15212 15026 15240 15302
rect 15200 15020 15252 15026
rect 15200 14962 15252 14968
rect 15384 14612 15436 14618
rect 15384 14554 15436 14560
rect 15016 14408 15068 14414
rect 15016 14350 15068 14356
rect 13452 13932 13504 13938
rect 13452 13874 13504 13880
rect 13268 13864 13320 13870
rect 13268 13806 13320 13812
rect 13176 12776 13228 12782
rect 13176 12718 13228 12724
rect 12624 11756 12676 11762
rect 12624 11698 12676 11704
rect 12900 11756 12952 11762
rect 12900 11698 12952 11704
rect 12256 11348 12308 11354
rect 12256 11290 12308 11296
rect 12268 10742 12296 11290
rect 12912 11218 12940 11698
rect 12900 11212 12952 11218
rect 12900 11154 12952 11160
rect 12256 10736 12308 10742
rect 12256 10678 12308 10684
rect 11796 10668 11848 10674
rect 11796 10610 11848 10616
rect 12164 10668 12216 10674
rect 12164 10610 12216 10616
rect 11612 10056 11664 10062
rect 11612 9998 11664 10004
rect 11336 9988 11388 9994
rect 11336 9930 11388 9936
rect 11348 9586 11376 9930
rect 11520 9920 11572 9926
rect 11520 9862 11572 9868
rect 11336 9580 11388 9586
rect 11336 9522 11388 9528
rect 11428 9580 11480 9586
rect 11428 9522 11480 9528
rect 11440 8090 11468 9522
rect 11532 9382 11560 9862
rect 11624 9518 11652 9998
rect 11808 9722 11836 10610
rect 12256 10124 12308 10130
rect 12256 10066 12308 10072
rect 11796 9716 11848 9722
rect 11796 9658 11848 9664
rect 12268 9586 12296 10066
rect 12912 10062 12940 11154
rect 13188 10674 13216 12718
rect 13280 12646 13308 13806
rect 13464 13326 13492 13874
rect 14924 13728 14976 13734
rect 14924 13670 14976 13676
rect 14556 13388 14608 13394
rect 14556 13330 14608 13336
rect 13452 13320 13504 13326
rect 13452 13262 13504 13268
rect 13268 12640 13320 12646
rect 13268 12582 13320 12588
rect 13464 12238 13492 13262
rect 14568 13258 14596 13330
rect 14936 13326 14964 13670
rect 15028 13376 15056 14350
rect 15292 14340 15344 14346
rect 15292 14282 15344 14288
rect 15108 13932 15160 13938
rect 15160 13892 15240 13920
rect 15108 13874 15160 13880
rect 15108 13388 15160 13394
rect 15028 13348 15108 13376
rect 14740 13320 14792 13326
rect 14738 13288 14740 13297
rect 14924 13320 14976 13326
rect 14792 13288 14794 13297
rect 14556 13252 14608 13258
rect 14924 13262 14976 13268
rect 14738 13223 14794 13232
rect 14556 13194 14608 13200
rect 14568 12782 14596 13194
rect 14740 12844 14792 12850
rect 14740 12786 14792 12792
rect 14556 12776 14608 12782
rect 14556 12718 14608 12724
rect 14752 12646 14780 12786
rect 14556 12640 14608 12646
rect 14556 12582 14608 12588
rect 14740 12640 14792 12646
rect 14740 12582 14792 12588
rect 13452 12232 13504 12238
rect 13452 12174 13504 12180
rect 13464 11762 13492 12174
rect 14568 12170 14596 12582
rect 14752 12442 14780 12582
rect 14740 12436 14792 12442
rect 14740 12378 14792 12384
rect 14752 12306 14780 12378
rect 14740 12300 14792 12306
rect 14740 12242 14792 12248
rect 14648 12232 14700 12238
rect 14648 12174 14700 12180
rect 14556 12164 14608 12170
rect 14556 12106 14608 12112
rect 14280 12096 14332 12102
rect 14280 12038 14332 12044
rect 14292 11762 14320 12038
rect 13452 11756 13504 11762
rect 13452 11698 13504 11704
rect 14280 11756 14332 11762
rect 14280 11698 14332 11704
rect 13464 11150 13492 11698
rect 14660 11694 14688 12174
rect 14740 12096 14792 12102
rect 14740 12038 14792 12044
rect 14648 11688 14700 11694
rect 14648 11630 14700 11636
rect 14752 11354 14780 12038
rect 14832 11756 14884 11762
rect 15028 11744 15056 13348
rect 15108 13330 15160 13336
rect 15108 13184 15160 13190
rect 15212 13172 15240 13892
rect 15304 13462 15332 14282
rect 15396 14006 15424 14554
rect 15568 14408 15620 14414
rect 15568 14350 15620 14356
rect 15384 14000 15436 14006
rect 15384 13942 15436 13948
rect 15384 13864 15436 13870
rect 15436 13824 15516 13852
rect 15384 13806 15436 13812
rect 15292 13456 15344 13462
rect 15292 13398 15344 13404
rect 15212 13144 15424 13172
rect 15108 13126 15160 13132
rect 15120 12866 15148 13126
rect 15120 12838 15332 12866
rect 15304 12442 15332 12838
rect 15292 12436 15344 12442
rect 15292 12378 15344 12384
rect 15200 12368 15252 12374
rect 15200 12310 15252 12316
rect 14884 11716 15148 11744
rect 14832 11698 14884 11704
rect 14740 11348 14792 11354
rect 14740 11290 14792 11296
rect 13452 11144 13504 11150
rect 13452 11086 13504 11092
rect 14280 11144 14332 11150
rect 14280 11086 14332 11092
rect 14372 11144 14424 11150
rect 14372 11086 14424 11092
rect 14096 11008 14148 11014
rect 14096 10950 14148 10956
rect 13176 10668 13228 10674
rect 13176 10610 13228 10616
rect 12900 10056 12952 10062
rect 12900 9998 12952 10004
rect 12348 9920 12400 9926
rect 12348 9862 12400 9868
rect 12256 9580 12308 9586
rect 12256 9522 12308 9528
rect 11612 9512 11664 9518
rect 11612 9454 11664 9460
rect 11520 9376 11572 9382
rect 11520 9318 11572 9324
rect 11624 8922 11652 9454
rect 12256 9036 12308 9042
rect 12256 8978 12308 8984
rect 11532 8894 11652 8922
rect 11532 8634 11560 8894
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 11428 8084 11480 8090
rect 11428 8026 11480 8032
rect 11336 7948 11388 7954
rect 11336 7890 11388 7896
rect 11348 6798 11376 7890
rect 11532 7886 11560 8570
rect 11612 8492 11664 8498
rect 11612 8434 11664 8440
rect 11980 8492 12032 8498
rect 11980 8434 12032 8440
rect 11624 8090 11652 8434
rect 11992 8090 12020 8434
rect 12268 8090 12296 8978
rect 12360 8974 12388 9862
rect 13188 9674 13216 10610
rect 14108 10606 14136 10950
rect 14096 10600 14148 10606
rect 14096 10542 14148 10548
rect 14188 10464 14240 10470
rect 14188 10406 14240 10412
rect 14200 10062 14228 10406
rect 14292 10146 14320 11086
rect 14384 10470 14412 11086
rect 15016 11008 15068 11014
rect 15016 10950 15068 10956
rect 15028 10742 15056 10950
rect 15016 10736 15068 10742
rect 15016 10678 15068 10684
rect 14832 10668 14884 10674
rect 14832 10610 14884 10616
rect 14740 10600 14792 10606
rect 14740 10542 14792 10548
rect 14372 10464 14424 10470
rect 14372 10406 14424 10412
rect 14292 10118 14412 10146
rect 14384 10062 14412 10118
rect 14188 10056 14240 10062
rect 14188 9998 14240 10004
rect 14372 10056 14424 10062
rect 14372 9998 14424 10004
rect 13096 9646 13216 9674
rect 13096 9586 13124 9646
rect 13084 9580 13136 9586
rect 13084 9522 13136 9528
rect 14752 9382 14780 10542
rect 14844 10266 14872 10610
rect 14832 10260 14884 10266
rect 14832 10202 14884 10208
rect 14740 9376 14792 9382
rect 14740 9318 14792 9324
rect 12348 8968 12400 8974
rect 12348 8910 12400 8916
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 13728 8968 13780 8974
rect 13728 8910 13780 8916
rect 12532 8832 12584 8838
rect 12532 8774 12584 8780
rect 11612 8084 11664 8090
rect 11612 8026 11664 8032
rect 11980 8084 12032 8090
rect 11980 8026 12032 8032
rect 12256 8084 12308 8090
rect 12256 8026 12308 8032
rect 12544 7886 12572 8774
rect 13556 8634 13584 8910
rect 13544 8628 13596 8634
rect 13544 8570 13596 8576
rect 13740 8566 13768 8910
rect 14752 8566 14780 9318
rect 15028 9178 15056 10678
rect 15120 10198 15148 11716
rect 15108 10192 15160 10198
rect 15108 10134 15160 10140
rect 15212 10130 15240 12310
rect 15396 10810 15424 13144
rect 15488 12986 15516 13824
rect 15476 12980 15528 12986
rect 15476 12922 15528 12928
rect 15476 12844 15528 12850
rect 15476 12786 15528 12792
rect 15488 12170 15516 12786
rect 15580 12646 15608 14350
rect 15752 13728 15804 13734
rect 15752 13670 15804 13676
rect 15764 13326 15792 13670
rect 15752 13320 15804 13326
rect 15750 13288 15752 13297
rect 15804 13288 15806 13297
rect 15750 13223 15806 13232
rect 15660 13184 15712 13190
rect 15660 13126 15712 13132
rect 15672 12782 15700 13126
rect 15660 12776 15712 12782
rect 15660 12718 15712 12724
rect 15568 12640 15620 12646
rect 15568 12582 15620 12588
rect 15476 12164 15528 12170
rect 15476 12106 15528 12112
rect 15476 11552 15528 11558
rect 15476 11494 15528 11500
rect 15488 11082 15516 11494
rect 15476 11076 15528 11082
rect 15476 11018 15528 11024
rect 15384 10804 15436 10810
rect 15384 10746 15436 10752
rect 15488 10674 15516 11018
rect 15856 10674 15884 17682
rect 16224 17338 16252 17682
rect 16212 17332 16264 17338
rect 16212 17274 16264 17280
rect 16500 16250 16528 18226
rect 16776 18154 16804 18634
rect 16764 18148 16816 18154
rect 16764 18090 16816 18096
rect 16868 17270 16896 20198
rect 16948 19372 17000 19378
rect 16948 19314 17000 19320
rect 16960 18834 16988 19314
rect 16948 18828 17000 18834
rect 16948 18770 17000 18776
rect 16960 18426 16988 18770
rect 16948 18420 17000 18426
rect 16948 18362 17000 18368
rect 17052 18358 17080 21814
rect 17316 21548 17368 21554
rect 17316 21490 17368 21496
rect 17328 21010 17356 21490
rect 17316 21004 17368 21010
rect 17316 20946 17368 20952
rect 17328 20602 17356 20946
rect 17316 20596 17368 20602
rect 17316 20538 17368 20544
rect 17132 20460 17184 20466
rect 17132 20402 17184 20408
rect 17144 19514 17172 20402
rect 17512 19990 17540 24142
rect 17592 23520 17644 23526
rect 17592 23462 17644 23468
rect 17604 23118 17632 23462
rect 17788 23254 17816 24550
rect 17972 23866 18000 25230
rect 18052 24812 18104 24818
rect 18052 24754 18104 24760
rect 17960 23860 18012 23866
rect 17960 23802 18012 23808
rect 18064 23474 18092 24754
rect 18156 24682 18184 25910
rect 18340 25702 18368 26794
rect 18524 26042 18552 27270
rect 18708 27033 18736 27814
rect 19720 27674 19748 27950
rect 19708 27668 19760 27674
rect 19708 27610 19760 27616
rect 19340 27532 19392 27538
rect 19340 27474 19392 27480
rect 19248 27396 19300 27402
rect 19248 27338 19300 27344
rect 18694 27024 18750 27033
rect 19260 26994 19288 27338
rect 18694 26959 18750 26968
rect 19248 26988 19300 26994
rect 19248 26930 19300 26936
rect 18512 26036 18564 26042
rect 18512 25978 18564 25984
rect 19260 25974 19288 26930
rect 19352 26518 19380 27474
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 19524 26920 19576 26926
rect 19522 26888 19524 26897
rect 19576 26888 19578 26897
rect 19996 26858 20024 28018
rect 20180 27606 20208 28478
rect 20260 28008 20312 28014
rect 20260 27950 20312 27956
rect 20168 27600 20220 27606
rect 20168 27542 20220 27548
rect 20168 27464 20220 27470
rect 20166 27432 20168 27441
rect 20220 27432 20222 27441
rect 20166 27367 20222 27376
rect 20168 27328 20220 27334
rect 20272 27316 20300 27950
rect 20364 27674 20392 29106
rect 20456 28694 20484 30631
rect 20536 28960 20588 28966
rect 20536 28902 20588 28908
rect 20444 28688 20496 28694
rect 20444 28630 20496 28636
rect 20444 28552 20496 28558
rect 20444 28494 20496 28500
rect 20352 27668 20404 27674
rect 20352 27610 20404 27616
rect 20220 27288 20300 27316
rect 20168 27270 20220 27276
rect 20076 26988 20128 26994
rect 20076 26930 20128 26936
rect 19522 26823 19578 26832
rect 19984 26852 20036 26858
rect 19984 26794 20036 26800
rect 19892 26784 19944 26790
rect 19892 26726 19944 26732
rect 19340 26512 19392 26518
rect 19340 26454 19392 26460
rect 19904 26382 19932 26726
rect 19892 26376 19944 26382
rect 19944 26324 20024 26330
rect 19892 26318 20024 26324
rect 19904 26302 20024 26318
rect 20088 26314 20116 26930
rect 20180 26761 20208 27270
rect 20364 27130 20392 27610
rect 20456 27169 20484 28494
rect 20548 27334 20576 28902
rect 20640 28558 20668 31726
rect 20720 31680 20772 31686
rect 20720 31622 20772 31628
rect 20732 31210 20760 31622
rect 21100 31278 21128 31758
rect 21824 31680 21876 31686
rect 21824 31622 21876 31628
rect 21916 31680 21968 31686
rect 21916 31622 21968 31628
rect 21836 31346 21864 31622
rect 21180 31340 21232 31346
rect 21180 31282 21232 31288
rect 21824 31340 21876 31346
rect 21824 31282 21876 31288
rect 21088 31272 21140 31278
rect 21088 31214 21140 31220
rect 20720 31204 20772 31210
rect 20720 31146 20772 31152
rect 21100 30938 21128 31214
rect 21088 30932 21140 30938
rect 21088 30874 21140 30880
rect 20812 30320 20864 30326
rect 20812 30262 20864 30268
rect 20720 29028 20772 29034
rect 20720 28970 20772 28976
rect 20732 28558 20760 28970
rect 20628 28552 20680 28558
rect 20628 28494 20680 28500
rect 20720 28552 20772 28558
rect 20720 28494 20772 28500
rect 20824 28370 20852 30262
rect 21192 29730 21220 31282
rect 21456 31204 21508 31210
rect 21456 31146 21508 31152
rect 21468 30734 21496 31146
rect 21456 30728 21508 30734
rect 21456 30670 21508 30676
rect 21272 30660 21324 30666
rect 21272 30602 21324 30608
rect 21284 29850 21312 30602
rect 21468 30394 21496 30670
rect 21640 30592 21692 30598
rect 21640 30534 21692 30540
rect 21732 30592 21784 30598
rect 21732 30534 21784 30540
rect 21456 30388 21508 30394
rect 21456 30330 21508 30336
rect 21652 30326 21680 30534
rect 21640 30320 21692 30326
rect 21640 30262 21692 30268
rect 21364 30252 21416 30258
rect 21364 30194 21416 30200
rect 21272 29844 21324 29850
rect 21272 29786 21324 29792
rect 21100 29702 21220 29730
rect 21100 29646 21128 29702
rect 21088 29640 21140 29646
rect 21088 29582 21140 29588
rect 21100 29238 21128 29582
rect 21088 29232 21140 29238
rect 21088 29174 21140 29180
rect 20904 29164 20956 29170
rect 20904 29106 20956 29112
rect 20916 28966 20944 29106
rect 20904 28960 20956 28966
rect 20904 28902 20956 28908
rect 20640 28342 20852 28370
rect 20640 28218 20668 28342
rect 20628 28212 20680 28218
rect 20628 28154 20680 28160
rect 20628 28076 20680 28082
rect 20628 28018 20680 28024
rect 20720 28076 20772 28082
rect 20916 28064 20944 28902
rect 21100 28234 21128 29174
rect 21100 28206 21312 28234
rect 21180 28076 21232 28082
rect 20772 28036 20944 28064
rect 20996 28042 21048 28048
rect 20720 28018 20772 28024
rect 20640 27538 20668 28018
rect 20628 27532 20680 27538
rect 20628 27474 20680 27480
rect 20732 27441 20760 28018
rect 20996 27984 21048 27990
rect 21100 28036 21180 28064
rect 21008 27674 21036 27984
rect 20996 27668 21048 27674
rect 20996 27610 21048 27616
rect 20718 27432 20774 27441
rect 20628 27396 20680 27402
rect 21100 27402 21128 28036
rect 21180 28018 21232 28024
rect 21284 28014 21312 28206
rect 21272 28008 21324 28014
rect 21272 27950 21324 27956
rect 20718 27367 20774 27376
rect 21088 27396 21140 27402
rect 20628 27338 20680 27344
rect 21088 27338 21140 27344
rect 20536 27328 20588 27334
rect 20536 27270 20588 27276
rect 20442 27160 20498 27169
rect 20260 27124 20312 27130
rect 20260 27066 20312 27072
rect 20352 27124 20404 27130
rect 20442 27095 20498 27104
rect 20352 27066 20404 27072
rect 20272 26926 20300 27066
rect 20640 26994 20668 27338
rect 20996 27056 21048 27062
rect 20996 26998 21048 27004
rect 20444 26988 20496 26994
rect 20444 26930 20496 26936
rect 20628 26988 20680 26994
rect 20628 26930 20680 26936
rect 20260 26920 20312 26926
rect 20260 26862 20312 26868
rect 20166 26752 20222 26761
rect 20166 26687 20222 26696
rect 20168 26376 20220 26382
rect 20168 26318 20220 26324
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 19248 25968 19300 25974
rect 19248 25910 19300 25916
rect 19996 25838 20024 26302
rect 20076 26308 20128 26314
rect 20076 26250 20128 26256
rect 20088 25906 20116 26250
rect 20180 25906 20208 26318
rect 20076 25900 20128 25906
rect 20076 25842 20128 25848
rect 20168 25900 20220 25906
rect 20168 25842 20220 25848
rect 19984 25832 20036 25838
rect 20456 25786 20484 26930
rect 21008 26382 21036 26998
rect 20720 26376 20772 26382
rect 20720 26318 20772 26324
rect 20996 26376 21048 26382
rect 20996 26318 21048 26324
rect 19984 25774 20036 25780
rect 20364 25770 20484 25786
rect 20352 25764 20484 25770
rect 20404 25758 20484 25764
rect 20352 25706 20404 25712
rect 18328 25696 18380 25702
rect 18328 25638 18380 25644
rect 19064 25696 19116 25702
rect 19064 25638 19116 25644
rect 18604 25152 18656 25158
rect 18604 25094 18656 25100
rect 18616 24818 18644 25094
rect 19076 24954 19104 25638
rect 19432 25288 19484 25294
rect 19432 25230 19484 25236
rect 20076 25288 20128 25294
rect 20076 25230 20128 25236
rect 18972 24948 19024 24954
rect 18972 24890 19024 24896
rect 19064 24948 19116 24954
rect 19064 24890 19116 24896
rect 18604 24812 18656 24818
rect 18604 24754 18656 24760
rect 18144 24676 18196 24682
rect 18144 24618 18196 24624
rect 18512 24200 18564 24206
rect 18512 24142 18564 24148
rect 18236 24064 18288 24070
rect 18236 24006 18288 24012
rect 18064 23446 18184 23474
rect 17776 23248 17828 23254
rect 17776 23190 17828 23196
rect 17592 23112 17644 23118
rect 17592 23054 17644 23060
rect 17960 23044 18012 23050
rect 17960 22986 18012 22992
rect 17684 22772 17736 22778
rect 17684 22714 17736 22720
rect 17696 21962 17724 22714
rect 17776 22228 17828 22234
rect 17776 22170 17828 22176
rect 17788 22030 17816 22170
rect 17776 22024 17828 22030
rect 17776 21966 17828 21972
rect 17684 21956 17736 21962
rect 17684 21898 17736 21904
rect 17788 20398 17816 21966
rect 17868 20528 17920 20534
rect 17868 20470 17920 20476
rect 17776 20392 17828 20398
rect 17776 20334 17828 20340
rect 17500 19984 17552 19990
rect 17500 19926 17552 19932
rect 17880 19922 17908 20470
rect 17868 19916 17920 19922
rect 17868 19858 17920 19864
rect 17972 19854 18000 22986
rect 18052 22500 18104 22506
rect 18052 22442 18104 22448
rect 18064 20466 18092 22442
rect 18156 21894 18184 23446
rect 18248 22030 18276 24006
rect 18524 22710 18552 24142
rect 18696 23792 18748 23798
rect 18696 23734 18748 23740
rect 18604 23656 18656 23662
rect 18604 23598 18656 23604
rect 18512 22704 18564 22710
rect 18512 22646 18564 22652
rect 18616 22642 18644 23598
rect 18604 22636 18656 22642
rect 18604 22578 18656 22584
rect 18236 22024 18288 22030
rect 18236 21966 18288 21972
rect 18144 21888 18196 21894
rect 18144 21830 18196 21836
rect 18326 21584 18382 21593
rect 18326 21519 18382 21528
rect 18602 21584 18658 21593
rect 18602 21519 18604 21528
rect 18052 20460 18104 20466
rect 18052 20402 18104 20408
rect 17960 19848 18012 19854
rect 17960 19790 18012 19796
rect 17132 19508 17184 19514
rect 17132 19450 17184 19456
rect 17144 18358 17172 19450
rect 17224 19372 17276 19378
rect 17224 19314 17276 19320
rect 17040 18352 17092 18358
rect 17040 18294 17092 18300
rect 17132 18352 17184 18358
rect 17132 18294 17184 18300
rect 17040 18216 17092 18222
rect 17040 18158 17092 18164
rect 16948 17604 17000 17610
rect 16948 17546 17000 17552
rect 16960 17270 16988 17546
rect 16856 17264 16908 17270
rect 16856 17206 16908 17212
rect 16948 17264 17000 17270
rect 16948 17206 17000 17212
rect 16960 16726 16988 17206
rect 17052 17202 17080 18158
rect 17236 18154 17264 19314
rect 17972 18902 18000 19790
rect 17960 18896 18012 18902
rect 17960 18838 18012 18844
rect 17960 18624 18012 18630
rect 17960 18566 18012 18572
rect 17224 18148 17276 18154
rect 17224 18090 17276 18096
rect 17868 17536 17920 17542
rect 17868 17478 17920 17484
rect 17132 17264 17184 17270
rect 17132 17206 17184 17212
rect 17040 17196 17092 17202
rect 17040 17138 17092 17144
rect 17052 17066 17080 17138
rect 17040 17060 17092 17066
rect 17040 17002 17092 17008
rect 16948 16720 17000 16726
rect 16948 16662 17000 16668
rect 16488 16244 16540 16250
rect 16488 16186 16540 16192
rect 16396 15972 16448 15978
rect 16396 15914 16448 15920
rect 16408 14618 16436 15914
rect 16672 15428 16724 15434
rect 16672 15370 16724 15376
rect 16684 15162 16712 15370
rect 16672 15156 16724 15162
rect 16672 15098 16724 15104
rect 16396 14612 16448 14618
rect 16396 14554 16448 14560
rect 16120 14272 16172 14278
rect 16120 14214 16172 14220
rect 16132 13938 16160 14214
rect 17144 13938 17172 17206
rect 17224 16992 17276 16998
rect 17224 16934 17276 16940
rect 17236 16590 17264 16934
rect 17880 16590 17908 17478
rect 17224 16584 17276 16590
rect 17224 16526 17276 16532
rect 17868 16584 17920 16590
rect 17868 16526 17920 16532
rect 17592 15904 17644 15910
rect 17592 15846 17644 15852
rect 17604 15026 17632 15846
rect 17972 15502 18000 18566
rect 18064 17678 18092 20402
rect 18236 19916 18288 19922
rect 18236 19858 18288 19864
rect 18248 18766 18276 19858
rect 18236 18760 18288 18766
rect 18236 18702 18288 18708
rect 18144 18692 18196 18698
rect 18144 18634 18196 18640
rect 18156 18426 18184 18634
rect 18144 18420 18196 18426
rect 18144 18362 18196 18368
rect 18248 18290 18276 18702
rect 18236 18284 18288 18290
rect 18236 18226 18288 18232
rect 18236 18080 18288 18086
rect 18236 18022 18288 18028
rect 18052 17672 18104 17678
rect 18104 17632 18184 17660
rect 18052 17614 18104 17620
rect 18156 16998 18184 17632
rect 18144 16992 18196 16998
rect 18144 16934 18196 16940
rect 18248 16726 18276 18022
rect 18340 17610 18368 21519
rect 18656 21519 18658 21528
rect 18604 21490 18656 21496
rect 18708 20534 18736 23734
rect 18984 23662 19012 24890
rect 19444 24682 19472 25230
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 19800 24812 19852 24818
rect 19800 24754 19852 24760
rect 19432 24676 19484 24682
rect 19432 24618 19484 24624
rect 19444 24410 19472 24618
rect 19812 24410 19840 24754
rect 19432 24404 19484 24410
rect 19432 24346 19484 24352
rect 19800 24404 19852 24410
rect 19800 24346 19852 24352
rect 19432 24064 19484 24070
rect 19432 24006 19484 24012
rect 19444 23730 19472 24006
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 19432 23724 19484 23730
rect 19432 23666 19484 23672
rect 18972 23656 19024 23662
rect 18972 23598 19024 23604
rect 19984 23588 20036 23594
rect 19984 23530 20036 23536
rect 19340 23520 19392 23526
rect 19340 23462 19392 23468
rect 18788 23316 18840 23322
rect 18788 23258 18840 23264
rect 18800 23118 18828 23258
rect 18788 23112 18840 23118
rect 18788 23054 18840 23060
rect 18696 20528 18748 20534
rect 18696 20470 18748 20476
rect 18708 18902 18736 20470
rect 18800 19378 18828 23054
rect 19064 22024 19116 22030
rect 19064 21966 19116 21972
rect 18880 21548 18932 21554
rect 18880 21490 18932 21496
rect 18788 19372 18840 19378
rect 18788 19314 18840 19320
rect 18696 18896 18748 18902
rect 18696 18838 18748 18844
rect 18420 18828 18472 18834
rect 18420 18770 18472 18776
rect 18432 18737 18460 18770
rect 18418 18728 18474 18737
rect 18418 18663 18474 18672
rect 18708 17814 18736 18838
rect 18696 17808 18748 17814
rect 18696 17750 18748 17756
rect 18328 17604 18380 17610
rect 18328 17546 18380 17552
rect 18340 17270 18368 17546
rect 18328 17264 18380 17270
rect 18328 17206 18380 17212
rect 18236 16720 18288 16726
rect 18236 16662 18288 16668
rect 18052 16040 18104 16046
rect 18052 15982 18104 15988
rect 17960 15496 18012 15502
rect 17960 15438 18012 15444
rect 17592 15020 17644 15026
rect 17592 14962 17644 14968
rect 17316 14408 17368 14414
rect 17316 14350 17368 14356
rect 16120 13932 16172 13938
rect 16120 13874 16172 13880
rect 17132 13932 17184 13938
rect 17132 13874 17184 13880
rect 16948 13252 17000 13258
rect 16948 13194 17000 13200
rect 16960 12850 16988 13194
rect 16948 12844 17000 12850
rect 16948 12786 17000 12792
rect 17328 12782 17356 14350
rect 18064 13938 18092 15982
rect 18248 15706 18276 16662
rect 18708 16590 18736 17750
rect 18696 16584 18748 16590
rect 18696 16526 18748 16532
rect 18696 16448 18748 16454
rect 18696 16390 18748 16396
rect 18708 16114 18736 16390
rect 18696 16108 18748 16114
rect 18696 16050 18748 16056
rect 18892 15978 18920 21490
rect 18972 20528 19024 20534
rect 18972 20470 19024 20476
rect 18984 18630 19012 20470
rect 18972 18624 19024 18630
rect 18972 18566 19024 18572
rect 19076 17542 19104 21966
rect 19352 21554 19380 23462
rect 19432 23112 19484 23118
rect 19432 23054 19484 23060
rect 19444 22778 19472 23054
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 19432 22772 19484 22778
rect 19432 22714 19484 22720
rect 19444 22030 19472 22714
rect 19432 22024 19484 22030
rect 19432 21966 19484 21972
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 19340 21548 19392 21554
rect 19340 21490 19392 21496
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 19432 20596 19484 20602
rect 19432 20538 19484 20544
rect 19340 19780 19392 19786
rect 19340 19722 19392 19728
rect 19248 19372 19300 19378
rect 19248 19314 19300 19320
rect 19156 19304 19208 19310
rect 19156 19246 19208 19252
rect 19168 18086 19196 19246
rect 19260 18290 19288 19314
rect 19352 18970 19380 19722
rect 19340 18964 19392 18970
rect 19340 18906 19392 18912
rect 19352 18358 19380 18906
rect 19340 18352 19392 18358
rect 19340 18294 19392 18300
rect 19248 18284 19300 18290
rect 19248 18226 19300 18232
rect 19156 18080 19208 18086
rect 19156 18022 19208 18028
rect 19064 17536 19116 17542
rect 19064 17478 19116 17484
rect 19168 17202 19196 18022
rect 19260 17626 19288 18226
rect 19260 17610 19380 17626
rect 19260 17604 19392 17610
rect 19260 17598 19340 17604
rect 19340 17546 19392 17552
rect 19156 17196 19208 17202
rect 19156 17138 19208 17144
rect 19168 16522 19196 17138
rect 19444 17082 19472 20538
rect 19996 19854 20024 23530
rect 20088 21690 20116 25230
rect 20168 24268 20220 24274
rect 20168 24210 20220 24216
rect 20076 21684 20128 21690
rect 20076 21626 20128 21632
rect 20180 21298 20208 24210
rect 20260 23180 20312 23186
rect 20260 23122 20312 23128
rect 20272 22642 20300 23122
rect 20260 22636 20312 22642
rect 20260 22578 20312 22584
rect 20260 22432 20312 22438
rect 20260 22374 20312 22380
rect 20272 22030 20300 22374
rect 20364 22098 20392 25706
rect 20732 25430 20760 26318
rect 20720 25424 20772 25430
rect 20720 25366 20772 25372
rect 21008 25294 21036 26318
rect 21100 25498 21128 27338
rect 21284 26450 21312 27950
rect 21272 26444 21324 26450
rect 21272 26386 21324 26392
rect 21376 26246 21404 30194
rect 21744 29102 21772 30534
rect 21836 30258 21864 31282
rect 21928 31210 21956 31622
rect 22008 31272 22060 31278
rect 22008 31214 22060 31220
rect 22744 31272 22796 31278
rect 22744 31214 22796 31220
rect 21916 31204 21968 31210
rect 21916 31146 21968 31152
rect 21824 30252 21876 30258
rect 21824 30194 21876 30200
rect 21928 29170 21956 31146
rect 22020 30258 22048 31214
rect 22192 30728 22244 30734
rect 22192 30670 22244 30676
rect 22376 30728 22428 30734
rect 22376 30670 22428 30676
rect 22100 30388 22152 30394
rect 22100 30330 22152 30336
rect 22008 30252 22060 30258
rect 22008 30194 22060 30200
rect 22112 29578 22140 30330
rect 22100 29572 22152 29578
rect 22100 29514 22152 29520
rect 21916 29164 21968 29170
rect 21916 29106 21968 29112
rect 21732 29096 21784 29102
rect 21732 29038 21784 29044
rect 21824 28552 21876 28558
rect 21824 28494 21876 28500
rect 22008 28552 22060 28558
rect 22008 28494 22060 28500
rect 21836 27878 21864 28494
rect 22020 28422 22048 28494
rect 22008 28416 22060 28422
rect 22008 28358 22060 28364
rect 21824 27872 21876 27878
rect 21824 27814 21876 27820
rect 21916 27464 21968 27470
rect 21916 27406 21968 27412
rect 21732 27396 21784 27402
rect 21732 27338 21784 27344
rect 21456 26444 21508 26450
rect 21456 26386 21508 26392
rect 21364 26240 21416 26246
rect 21364 26182 21416 26188
rect 21376 25906 21404 26182
rect 21468 26042 21496 26386
rect 21744 26246 21772 27338
rect 21928 26586 21956 27406
rect 22020 27062 22048 28358
rect 22112 28082 22140 29514
rect 22204 29306 22232 30670
rect 22192 29300 22244 29306
rect 22192 29242 22244 29248
rect 22388 28762 22416 30670
rect 22756 30394 22784 31214
rect 23032 30870 23060 32370
rect 23216 32026 23244 32710
rect 23676 32570 23704 32846
rect 23664 32564 23716 32570
rect 23664 32506 23716 32512
rect 23768 32450 23796 32914
rect 24124 32836 24176 32842
rect 24124 32778 24176 32784
rect 23572 32428 23624 32434
rect 23572 32370 23624 32376
rect 23676 32422 23796 32450
rect 23204 32020 23256 32026
rect 23204 31962 23256 31968
rect 23388 31680 23440 31686
rect 23388 31622 23440 31628
rect 23480 31680 23532 31686
rect 23480 31622 23532 31628
rect 23112 31340 23164 31346
rect 23112 31282 23164 31288
rect 23124 30938 23152 31282
rect 23204 31136 23256 31142
rect 23204 31078 23256 31084
rect 23112 30932 23164 30938
rect 23112 30874 23164 30880
rect 23020 30864 23072 30870
rect 23020 30806 23072 30812
rect 22836 30660 22888 30666
rect 22836 30602 22888 30608
rect 22744 30388 22796 30394
rect 22744 30330 22796 30336
rect 22744 30252 22796 30258
rect 22744 30194 22796 30200
rect 22468 30116 22520 30122
rect 22468 30058 22520 30064
rect 22480 29782 22508 30058
rect 22652 30048 22704 30054
rect 22652 29990 22704 29996
rect 22468 29776 22520 29782
rect 22468 29718 22520 29724
rect 22480 29510 22508 29718
rect 22468 29504 22520 29510
rect 22468 29446 22520 29452
rect 22376 28756 22428 28762
rect 22376 28698 22428 28704
rect 22100 28076 22152 28082
rect 22100 28018 22152 28024
rect 22008 27056 22060 27062
rect 22008 26998 22060 27004
rect 21916 26580 21968 26586
rect 21916 26522 21968 26528
rect 21916 26376 21968 26382
rect 21916 26318 21968 26324
rect 21732 26240 21784 26246
rect 21732 26182 21784 26188
rect 21456 26036 21508 26042
rect 21456 25978 21508 25984
rect 21364 25900 21416 25906
rect 21364 25842 21416 25848
rect 21928 25838 21956 26318
rect 21916 25832 21968 25838
rect 21916 25774 21968 25780
rect 21088 25492 21140 25498
rect 21088 25434 21140 25440
rect 21928 25362 21956 25774
rect 21916 25356 21968 25362
rect 21916 25298 21968 25304
rect 20996 25288 21048 25294
rect 20996 25230 21048 25236
rect 21364 25220 21416 25226
rect 21364 25162 21416 25168
rect 20534 24848 20590 24857
rect 20444 24812 20496 24818
rect 20534 24783 20536 24792
rect 20444 24754 20496 24760
rect 20588 24783 20590 24792
rect 21180 24812 21232 24818
rect 20536 24754 20588 24760
rect 21180 24754 21232 24760
rect 21272 24812 21324 24818
rect 21272 24754 21324 24760
rect 20456 24410 20484 24754
rect 20720 24608 20772 24614
rect 20720 24550 20772 24556
rect 20444 24404 20496 24410
rect 20444 24346 20496 24352
rect 20442 24304 20498 24313
rect 20442 24239 20444 24248
rect 20496 24239 20498 24248
rect 20444 24210 20496 24216
rect 20442 24168 20498 24177
rect 20732 24138 20760 24550
rect 20996 24200 21048 24206
rect 20996 24142 21048 24148
rect 20442 24103 20444 24112
rect 20496 24103 20498 24112
rect 20720 24132 20772 24138
rect 20444 24074 20496 24080
rect 20720 24074 20772 24080
rect 20444 23656 20496 23662
rect 20444 23598 20496 23604
rect 20352 22092 20404 22098
rect 20352 22034 20404 22040
rect 20260 22024 20312 22030
rect 20456 22001 20484 23598
rect 21008 23322 21036 24142
rect 21192 24041 21220 24754
rect 21284 24682 21312 24754
rect 21272 24676 21324 24682
rect 21272 24618 21324 24624
rect 21178 24032 21234 24041
rect 21178 23967 21234 23976
rect 21376 23866 21404 25162
rect 21732 24812 21784 24818
rect 21732 24754 21784 24760
rect 21364 23860 21416 23866
rect 21364 23802 21416 23808
rect 21088 23724 21140 23730
rect 21088 23666 21140 23672
rect 21100 23633 21128 23666
rect 21086 23624 21142 23633
rect 21086 23559 21142 23568
rect 21546 23352 21602 23361
rect 20996 23316 21048 23322
rect 21546 23287 21602 23296
rect 20996 23258 21048 23264
rect 21560 23118 21588 23287
rect 21744 23254 21772 24754
rect 21824 24608 21876 24614
rect 21822 24576 21824 24585
rect 21876 24576 21878 24585
rect 21822 24511 21878 24520
rect 21824 24200 21876 24206
rect 21824 24142 21876 24148
rect 21732 23248 21784 23254
rect 21732 23190 21784 23196
rect 20812 23112 20864 23118
rect 20812 23054 20864 23060
rect 21548 23112 21600 23118
rect 21548 23054 21600 23060
rect 20720 22636 20772 22642
rect 20720 22578 20772 22584
rect 20732 22234 20760 22578
rect 20720 22228 20772 22234
rect 20720 22170 20772 22176
rect 20260 21966 20312 21972
rect 20442 21992 20498 22001
rect 20442 21927 20498 21936
rect 20180 21270 20300 21298
rect 20076 20936 20128 20942
rect 20076 20878 20128 20884
rect 20088 20534 20116 20878
rect 20076 20528 20128 20534
rect 20076 20470 20128 20476
rect 20076 20052 20128 20058
rect 20076 19994 20128 20000
rect 19984 19848 20036 19854
rect 19984 19790 20036 19796
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 19984 19508 20036 19514
rect 19984 19450 20036 19456
rect 19800 19440 19852 19446
rect 19798 19408 19800 19417
rect 19852 19408 19854 19417
rect 19798 19343 19854 19352
rect 19800 19304 19852 19310
rect 19798 19272 19800 19281
rect 19852 19272 19854 19281
rect 19798 19207 19854 19216
rect 19706 18864 19762 18873
rect 19706 18799 19762 18808
rect 19720 18766 19748 18799
rect 19708 18760 19760 18766
rect 19708 18702 19760 18708
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 19524 17672 19576 17678
rect 19524 17614 19576 17620
rect 19536 17524 19564 17614
rect 19516 17496 19564 17524
rect 19516 17252 19544 17496
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 19516 17224 19564 17252
rect 19536 17134 19564 17224
rect 19352 17054 19472 17082
rect 19524 17128 19576 17134
rect 19524 17070 19576 17076
rect 19352 16674 19380 17054
rect 19432 16992 19484 16998
rect 19432 16934 19484 16940
rect 19260 16646 19380 16674
rect 19156 16516 19208 16522
rect 19156 16458 19208 16464
rect 19260 16130 19288 16646
rect 19340 16584 19392 16590
rect 19340 16526 19392 16532
rect 19352 16250 19380 16526
rect 19340 16244 19392 16250
rect 19340 16186 19392 16192
rect 19260 16114 19380 16130
rect 19260 16108 19392 16114
rect 19260 16102 19340 16108
rect 19340 16050 19392 16056
rect 19156 16040 19208 16046
rect 19156 15982 19208 15988
rect 18880 15972 18932 15978
rect 18880 15914 18932 15920
rect 18236 15700 18288 15706
rect 18236 15642 18288 15648
rect 18248 15094 18276 15642
rect 19168 15638 19196 15982
rect 19156 15632 19208 15638
rect 19156 15574 19208 15580
rect 19444 15502 19472 16934
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 19432 15496 19484 15502
rect 19432 15438 19484 15444
rect 18420 15360 18472 15366
rect 18420 15302 18472 15308
rect 18236 15088 18288 15094
rect 18236 15030 18288 15036
rect 18052 13932 18104 13938
rect 18104 13892 18184 13920
rect 18052 13874 18104 13880
rect 17960 13796 18012 13802
rect 17960 13738 18012 13744
rect 17972 13394 18000 13738
rect 18052 13728 18104 13734
rect 18052 13670 18104 13676
rect 17960 13388 18012 13394
rect 17960 13330 18012 13336
rect 17972 13190 18000 13330
rect 18064 13326 18092 13670
rect 18156 13394 18184 13892
rect 18144 13388 18196 13394
rect 18144 13330 18196 13336
rect 18052 13320 18104 13326
rect 18052 13262 18104 13268
rect 17960 13184 18012 13190
rect 17960 13126 18012 13132
rect 18144 12912 18196 12918
rect 18144 12854 18196 12860
rect 16764 12776 16816 12782
rect 16764 12718 16816 12724
rect 17316 12776 17368 12782
rect 17316 12718 17368 12724
rect 16488 12164 16540 12170
rect 16488 12106 16540 12112
rect 16500 11762 16528 12106
rect 16488 11756 16540 11762
rect 16488 11698 16540 11704
rect 16120 11688 16172 11694
rect 16120 11630 16172 11636
rect 16132 11150 16160 11630
rect 16672 11212 16724 11218
rect 16672 11154 16724 11160
rect 16120 11144 16172 11150
rect 16120 11086 16172 11092
rect 16580 11144 16632 11150
rect 16580 11086 16632 11092
rect 16132 10810 16160 11086
rect 16120 10804 16172 10810
rect 16120 10746 16172 10752
rect 15476 10668 15528 10674
rect 15476 10610 15528 10616
rect 15844 10668 15896 10674
rect 15844 10610 15896 10616
rect 15200 10124 15252 10130
rect 15200 10066 15252 10072
rect 15212 9500 15240 10066
rect 16592 9994 16620 11086
rect 16684 10266 16712 11154
rect 16776 11150 16804 12718
rect 17222 12472 17278 12481
rect 17222 12407 17224 12416
rect 17276 12407 17278 12416
rect 17224 12378 17276 12384
rect 16764 11144 16816 11150
rect 16764 11086 16816 11092
rect 16856 11076 16908 11082
rect 16856 11018 16908 11024
rect 16868 10810 16896 11018
rect 16856 10804 16908 10810
rect 16856 10746 16908 10752
rect 16672 10260 16724 10266
rect 16672 10202 16724 10208
rect 15384 9988 15436 9994
rect 15384 9930 15436 9936
rect 15936 9988 15988 9994
rect 15936 9930 15988 9936
rect 16580 9988 16632 9994
rect 16580 9930 16632 9936
rect 15396 9586 15424 9930
rect 15948 9722 15976 9930
rect 15936 9716 15988 9722
rect 15936 9658 15988 9664
rect 15384 9580 15436 9586
rect 15384 9522 15436 9528
rect 15292 9512 15344 9518
rect 15212 9472 15292 9500
rect 15292 9454 15344 9460
rect 16212 9512 16264 9518
rect 16212 9454 16264 9460
rect 15016 9172 15068 9178
rect 15016 9114 15068 9120
rect 13728 8560 13780 8566
rect 13728 8502 13780 8508
rect 14740 8560 14792 8566
rect 14740 8502 14792 8508
rect 13740 8430 13768 8502
rect 15304 8498 15332 9454
rect 16224 8974 16252 9454
rect 16212 8968 16264 8974
rect 16212 8910 16264 8916
rect 15292 8492 15344 8498
rect 15292 8434 15344 8440
rect 13728 8424 13780 8430
rect 13728 8366 13780 8372
rect 16592 8362 16620 9930
rect 16672 9512 16724 9518
rect 16672 9454 16724 9460
rect 16684 9110 16712 9454
rect 16672 9104 16724 9110
rect 16672 9046 16724 9052
rect 16684 8634 16712 9046
rect 16764 8832 16816 8838
rect 16764 8774 16816 8780
rect 16672 8628 16724 8634
rect 16672 8570 16724 8576
rect 16776 8566 16804 8774
rect 16764 8560 16816 8566
rect 16764 8502 16816 8508
rect 16580 8356 16632 8362
rect 16580 8298 16632 8304
rect 16592 7954 16620 8298
rect 17236 8090 17264 12378
rect 17328 12170 17356 12718
rect 17316 12164 17368 12170
rect 17316 12106 17368 12112
rect 18156 11286 18184 12854
rect 18432 12306 18460 15302
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 19996 15026 20024 19450
rect 20088 16794 20116 19994
rect 20168 19780 20220 19786
rect 20168 19722 20220 19728
rect 20180 19553 20208 19722
rect 20166 19544 20222 19553
rect 20166 19479 20222 19488
rect 20180 18986 20208 19479
rect 20272 19174 20300 21270
rect 20350 19544 20406 19553
rect 20350 19479 20352 19488
rect 20404 19479 20406 19488
rect 20352 19450 20404 19456
rect 20352 19304 20404 19310
rect 20352 19246 20404 19252
rect 20260 19168 20312 19174
rect 20260 19110 20312 19116
rect 20364 18986 20392 19246
rect 20180 18958 20392 18986
rect 20168 18284 20220 18290
rect 20168 18226 20220 18232
rect 20180 17882 20208 18226
rect 20168 17876 20220 17882
rect 20168 17818 20220 17824
rect 20456 17610 20484 21927
rect 20824 21894 20852 23054
rect 21836 22094 21864 24142
rect 22112 24138 22140 28018
rect 22388 27946 22416 28698
rect 22664 28558 22692 29990
rect 22756 29646 22784 30194
rect 22848 30054 22876 30602
rect 23124 30190 23152 30874
rect 23216 30802 23244 31078
rect 23204 30796 23256 30802
rect 23204 30738 23256 30744
rect 23204 30388 23256 30394
rect 23204 30330 23256 30336
rect 23112 30184 23164 30190
rect 23112 30126 23164 30132
rect 22836 30048 22888 30054
rect 22836 29990 22888 29996
rect 22928 30048 22980 30054
rect 22928 29990 22980 29996
rect 22836 29844 22888 29850
rect 22836 29786 22888 29792
rect 22744 29640 22796 29646
rect 22744 29582 22796 29588
rect 22848 28937 22876 29786
rect 22834 28928 22890 28937
rect 22834 28863 22890 28872
rect 22652 28552 22704 28558
rect 22652 28494 22704 28500
rect 22744 28076 22796 28082
rect 22744 28018 22796 28024
rect 22376 27940 22428 27946
rect 22376 27882 22428 27888
rect 22284 27872 22336 27878
rect 22284 27814 22336 27820
rect 22296 25838 22324 27814
rect 22560 27328 22612 27334
rect 22560 27270 22612 27276
rect 22374 27024 22430 27033
rect 22374 26959 22376 26968
rect 22428 26959 22430 26968
rect 22376 26930 22428 26936
rect 22468 26512 22520 26518
rect 22468 26454 22520 26460
rect 22376 25900 22428 25906
rect 22376 25842 22428 25848
rect 22284 25832 22336 25838
rect 22284 25774 22336 25780
rect 22190 24576 22246 24585
rect 22190 24511 22246 24520
rect 22204 24410 22232 24511
rect 22192 24404 22244 24410
rect 22192 24346 22244 24352
rect 22388 24274 22416 25842
rect 22376 24268 22428 24274
rect 22376 24210 22428 24216
rect 22100 24132 22152 24138
rect 22100 24074 22152 24080
rect 22098 23896 22154 23905
rect 22098 23831 22154 23840
rect 22112 23730 22140 23831
rect 22100 23724 22152 23730
rect 22100 23666 22152 23672
rect 22480 23662 22508 26454
rect 22572 25294 22600 27270
rect 22756 26926 22784 28018
rect 22744 26920 22796 26926
rect 22744 26862 22796 26868
rect 22652 25424 22704 25430
rect 22652 25366 22704 25372
rect 22560 25288 22612 25294
rect 22560 25230 22612 25236
rect 22560 24744 22612 24750
rect 22560 24686 22612 24692
rect 22572 23866 22600 24686
rect 22560 23860 22612 23866
rect 22560 23802 22612 23808
rect 22468 23656 22520 23662
rect 22466 23624 22468 23633
rect 22520 23624 22522 23633
rect 22466 23559 22522 23568
rect 22664 22778 22692 25366
rect 22848 25362 22876 28863
rect 22836 25356 22888 25362
rect 22836 25298 22888 25304
rect 22744 24608 22796 24614
rect 22742 24576 22744 24585
rect 22796 24576 22798 24585
rect 22742 24511 22798 24520
rect 22742 23896 22798 23905
rect 22742 23831 22798 23840
rect 22756 23730 22784 23831
rect 22744 23724 22796 23730
rect 22744 23666 22796 23672
rect 22744 23044 22796 23050
rect 22744 22986 22796 22992
rect 22652 22772 22704 22778
rect 22652 22714 22704 22720
rect 22756 22642 22784 22986
rect 22744 22636 22796 22642
rect 22744 22578 22796 22584
rect 22192 22500 22244 22506
rect 22192 22442 22244 22448
rect 22008 22432 22060 22438
rect 22008 22374 22060 22380
rect 22100 22432 22152 22438
rect 22100 22374 22152 22380
rect 21836 22066 21956 22094
rect 21548 21956 21600 21962
rect 21548 21898 21600 21904
rect 20812 21888 20864 21894
rect 20812 21830 20864 21836
rect 21560 21842 21588 21898
rect 21824 21888 21876 21894
rect 21560 21814 21680 21842
rect 21824 21830 21876 21836
rect 20812 21344 20864 21350
rect 20812 21286 20864 21292
rect 20720 20800 20772 20806
rect 20720 20742 20772 20748
rect 20732 20534 20760 20742
rect 20720 20528 20772 20534
rect 20720 20470 20772 20476
rect 20824 20466 20852 21286
rect 21652 21010 21680 21814
rect 21836 21554 21864 21830
rect 21824 21548 21876 21554
rect 21824 21490 21876 21496
rect 21640 21004 21692 21010
rect 21640 20946 21692 20952
rect 20904 20800 20956 20806
rect 20904 20742 20956 20748
rect 20812 20460 20864 20466
rect 20812 20402 20864 20408
rect 20628 20324 20680 20330
rect 20628 20266 20680 20272
rect 20640 19854 20668 20266
rect 20628 19848 20680 19854
rect 20628 19790 20680 19796
rect 20536 19712 20588 19718
rect 20536 19654 20588 19660
rect 20548 19378 20576 19654
rect 20916 19446 20944 20742
rect 20996 20596 21048 20602
rect 20996 20538 21048 20544
rect 21008 19922 21036 20538
rect 21180 20528 21232 20534
rect 21180 20470 21232 20476
rect 20996 19916 21048 19922
rect 20996 19858 21048 19864
rect 20904 19440 20956 19446
rect 20904 19382 20956 19388
rect 20536 19372 20588 19378
rect 20536 19314 20588 19320
rect 20534 19272 20590 19281
rect 21008 19242 21036 19858
rect 21192 19854 21220 20470
rect 21180 19848 21232 19854
rect 21180 19790 21232 19796
rect 21088 19508 21140 19514
rect 21088 19450 21140 19456
rect 20534 19207 20536 19216
rect 20588 19207 20590 19216
rect 20996 19236 21048 19242
rect 20536 19178 20588 19184
rect 20996 19178 21048 19184
rect 20812 19168 20864 19174
rect 20812 19110 20864 19116
rect 20824 17678 20852 19110
rect 20904 18828 20956 18834
rect 20904 18770 20956 18776
rect 20812 17672 20864 17678
rect 20812 17614 20864 17620
rect 20444 17604 20496 17610
rect 20444 17546 20496 17552
rect 20168 17536 20220 17542
rect 20168 17478 20220 17484
rect 20180 17202 20208 17478
rect 20916 17202 20944 18770
rect 20168 17196 20220 17202
rect 20168 17138 20220 17144
rect 20904 17196 20956 17202
rect 20904 17138 20956 17144
rect 20260 16992 20312 16998
rect 20260 16934 20312 16940
rect 20076 16788 20128 16794
rect 20076 16730 20128 16736
rect 20272 16114 20300 16934
rect 20260 16108 20312 16114
rect 20260 16050 20312 16056
rect 20260 15360 20312 15366
rect 20260 15302 20312 15308
rect 20812 15360 20864 15366
rect 20812 15302 20864 15308
rect 19984 15020 20036 15026
rect 19984 14962 20036 14968
rect 19156 14952 19208 14958
rect 19156 14894 19208 14900
rect 18972 14816 19024 14822
rect 18972 14758 19024 14764
rect 18880 14612 18932 14618
rect 18880 14554 18932 14560
rect 18892 14006 18920 14554
rect 18984 14074 19012 14758
rect 18972 14068 19024 14074
rect 18972 14010 19024 14016
rect 18880 14000 18932 14006
rect 18880 13942 18932 13948
rect 18604 13796 18656 13802
rect 18604 13738 18656 13744
rect 18616 12782 18644 13738
rect 19168 13172 19196 14894
rect 19432 14408 19484 14414
rect 19432 14350 19484 14356
rect 19340 14272 19392 14278
rect 19260 14232 19340 14260
rect 19260 13394 19288 14232
rect 19340 14214 19392 14220
rect 19444 13462 19472 14350
rect 19984 14340 20036 14346
rect 19984 14282 20036 14288
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 19996 14074 20024 14282
rect 19984 14068 20036 14074
rect 19984 14010 20036 14016
rect 19432 13456 19484 13462
rect 19432 13398 19484 13404
rect 19248 13388 19300 13394
rect 19248 13330 19300 13336
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 19248 13184 19300 13190
rect 19168 13144 19248 13172
rect 19248 13126 19300 13132
rect 18604 12776 18656 12782
rect 18604 12718 18656 12724
rect 18616 12306 18644 12718
rect 18696 12640 18748 12646
rect 18696 12582 18748 12588
rect 18708 12306 18736 12582
rect 18420 12300 18472 12306
rect 18420 12242 18472 12248
rect 18604 12300 18656 12306
rect 18604 12242 18656 12248
rect 18696 12300 18748 12306
rect 18696 12242 18748 12248
rect 19260 11694 19288 13126
rect 19340 12640 19392 12646
rect 19340 12582 19392 12588
rect 19352 11762 19380 12582
rect 19444 12442 19472 13262
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 20272 12986 20300 15302
rect 20352 15020 20404 15026
rect 20352 14962 20404 14968
rect 20364 14074 20392 14962
rect 20444 14816 20496 14822
rect 20444 14758 20496 14764
rect 20352 14068 20404 14074
rect 20352 14010 20404 14016
rect 20456 13938 20484 14758
rect 20824 14006 20852 15302
rect 20812 14000 20864 14006
rect 20812 13942 20864 13948
rect 20444 13932 20496 13938
rect 20444 13874 20496 13880
rect 20260 12980 20312 12986
rect 20260 12922 20312 12928
rect 20916 12918 20944 17138
rect 20996 16720 21048 16726
rect 20996 16662 21048 16668
rect 21008 15094 21036 16662
rect 21100 15502 21128 19450
rect 21456 17672 21508 17678
rect 21456 17614 21508 17620
rect 21468 17134 21496 17614
rect 21456 17128 21508 17134
rect 21456 17070 21508 17076
rect 21468 16590 21496 17070
rect 21456 16584 21508 16590
rect 21456 16526 21508 16532
rect 21468 15706 21496 16526
rect 21456 15700 21508 15706
rect 21456 15642 21508 15648
rect 21088 15496 21140 15502
rect 21088 15438 21140 15444
rect 20996 15088 21048 15094
rect 20996 15030 21048 15036
rect 21088 14816 21140 14822
rect 21088 14758 21140 14764
rect 21364 14816 21416 14822
rect 21364 14758 21416 14764
rect 21100 13870 21128 14758
rect 21376 14414 21404 14758
rect 21364 14408 21416 14414
rect 21364 14350 21416 14356
rect 21088 13864 21140 13870
rect 21088 13806 21140 13812
rect 21376 13326 21404 14350
rect 21456 14272 21508 14278
rect 21456 14214 21508 14220
rect 21468 14074 21496 14214
rect 21456 14068 21508 14074
rect 21456 14010 21508 14016
rect 21088 13320 21140 13326
rect 21088 13262 21140 13268
rect 21364 13320 21416 13326
rect 21364 13262 21416 13268
rect 20904 12912 20956 12918
rect 20904 12854 20956 12860
rect 20628 12844 20680 12850
rect 20628 12786 20680 12792
rect 20640 12442 20668 12786
rect 19432 12436 19484 12442
rect 19432 12378 19484 12384
rect 20628 12436 20680 12442
rect 20628 12378 20680 12384
rect 21100 12186 21128 13262
rect 21008 12158 21128 12186
rect 21364 12232 21416 12238
rect 21364 12174 21416 12180
rect 21008 12102 21036 12158
rect 20720 12096 20772 12102
rect 20720 12038 20772 12044
rect 20996 12096 21048 12102
rect 20996 12038 21048 12044
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 19340 11756 19392 11762
rect 19340 11698 19392 11704
rect 19248 11688 19300 11694
rect 19248 11630 19300 11636
rect 18144 11280 18196 11286
rect 18144 11222 18196 11228
rect 18512 11280 18564 11286
rect 18512 11222 18564 11228
rect 19340 11280 19392 11286
rect 19340 11222 19392 11228
rect 18236 11008 18288 11014
rect 18236 10950 18288 10956
rect 17960 10736 18012 10742
rect 18248 10690 18276 10950
rect 18012 10684 18276 10690
rect 17960 10678 18276 10684
rect 18420 10736 18472 10742
rect 18420 10678 18472 10684
rect 17972 10674 18276 10678
rect 17972 10668 18288 10674
rect 17972 10662 18236 10668
rect 18236 10610 18288 10616
rect 18144 10600 18196 10606
rect 18144 10542 18196 10548
rect 17960 10464 18012 10470
rect 17960 10406 18012 10412
rect 17972 10266 18000 10406
rect 17960 10260 18012 10266
rect 17960 10202 18012 10208
rect 18052 10192 18104 10198
rect 18052 10134 18104 10140
rect 17776 10056 17828 10062
rect 17776 9998 17828 10004
rect 17788 9110 17816 9998
rect 17776 9104 17828 9110
rect 17776 9046 17828 9052
rect 18064 8906 18092 10134
rect 18156 9178 18184 10542
rect 18432 9926 18460 10678
rect 18524 10606 18552 11222
rect 18604 11144 18656 11150
rect 18604 11086 18656 11092
rect 18512 10600 18564 10606
rect 18512 10542 18564 10548
rect 18616 10062 18644 11086
rect 19064 10124 19116 10130
rect 19064 10066 19116 10072
rect 18604 10056 18656 10062
rect 18604 9998 18656 10004
rect 18420 9920 18472 9926
rect 18420 9862 18472 9868
rect 18432 9654 18460 9862
rect 18420 9648 18472 9654
rect 18420 9590 18472 9596
rect 19076 9450 19104 10066
rect 19352 10062 19380 11222
rect 20732 11218 20760 12038
rect 21376 11898 21404 12174
rect 21364 11892 21416 11898
rect 21364 11834 21416 11840
rect 20812 11552 20864 11558
rect 20812 11494 20864 11500
rect 20720 11212 20772 11218
rect 20720 11154 20772 11160
rect 19432 11144 19484 11150
rect 19432 11086 19484 11092
rect 19248 10056 19300 10062
rect 19248 9998 19300 10004
rect 19340 10056 19392 10062
rect 19340 9998 19392 10004
rect 19260 9654 19288 9998
rect 19248 9648 19300 9654
rect 19248 9590 19300 9596
rect 19064 9444 19116 9450
rect 19064 9386 19116 9392
rect 18144 9172 18196 9178
rect 18144 9114 18196 9120
rect 19076 8974 19104 9386
rect 19444 9178 19472 11086
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 19984 10804 20036 10810
rect 19984 10746 20036 10752
rect 19892 10600 19944 10606
rect 19996 10588 20024 10746
rect 20168 10668 20220 10674
rect 20168 10610 20220 10616
rect 19944 10560 20024 10588
rect 19892 10542 19944 10548
rect 20180 10470 20208 10610
rect 20168 10464 20220 10470
rect 20168 10406 20220 10412
rect 20180 10266 20208 10406
rect 20168 10260 20220 10266
rect 20168 10202 20220 10208
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 19432 9172 19484 9178
rect 19432 9114 19484 9120
rect 20180 9042 20208 10202
rect 20732 10130 20760 11154
rect 20824 11150 20852 11494
rect 20812 11144 20864 11150
rect 20812 11086 20864 11092
rect 21652 11014 21680 20946
rect 21732 20936 21784 20942
rect 21732 20878 21784 20884
rect 21744 20602 21772 20878
rect 21928 20602 21956 22066
rect 22020 21962 22048 22374
rect 22008 21956 22060 21962
rect 22008 21898 22060 21904
rect 22112 21842 22140 22374
rect 22020 21814 22140 21842
rect 22020 21593 22048 21814
rect 22204 21622 22232 22442
rect 22652 22432 22704 22438
rect 22652 22374 22704 22380
rect 22664 22234 22692 22374
rect 22756 22234 22784 22578
rect 22652 22228 22704 22234
rect 22652 22170 22704 22176
rect 22744 22228 22796 22234
rect 22744 22170 22796 22176
rect 22192 21616 22244 21622
rect 22006 21584 22062 21593
rect 22192 21558 22244 21564
rect 22006 21519 22062 21528
rect 21732 20596 21784 20602
rect 21732 20538 21784 20544
rect 21916 20596 21968 20602
rect 21916 20538 21968 20544
rect 22020 20466 22048 21519
rect 22204 21078 22232 21558
rect 22560 21548 22612 21554
rect 22560 21490 22612 21496
rect 22284 21344 22336 21350
rect 22284 21286 22336 21292
rect 22192 21072 22244 21078
rect 22112 21020 22192 21026
rect 22112 21014 22244 21020
rect 22112 20998 22232 21014
rect 22112 20466 22140 20998
rect 22192 20528 22244 20534
rect 22192 20470 22244 20476
rect 22008 20460 22060 20466
rect 22008 20402 22060 20408
rect 22100 20460 22152 20466
rect 22100 20402 22152 20408
rect 22100 20052 22152 20058
rect 22100 19994 22152 20000
rect 21916 19304 21968 19310
rect 21916 19246 21968 19252
rect 21928 18766 21956 19246
rect 22008 18964 22060 18970
rect 22008 18906 22060 18912
rect 21916 18760 21968 18766
rect 21916 18702 21968 18708
rect 21928 18630 21956 18702
rect 21824 18624 21876 18630
rect 21824 18566 21876 18572
rect 21916 18624 21968 18630
rect 21916 18566 21968 18572
rect 21836 18290 21864 18566
rect 21824 18284 21876 18290
rect 21824 18226 21876 18232
rect 21928 18204 21956 18566
rect 22020 18290 22048 18906
rect 22008 18284 22060 18290
rect 22008 18226 22060 18232
rect 21919 18176 21956 18204
rect 21919 18170 21947 18176
rect 21836 18142 21947 18170
rect 21836 17882 21864 18142
rect 21824 17876 21876 17882
rect 21824 17818 21876 17824
rect 21916 17876 21968 17882
rect 21916 17818 21968 17824
rect 21822 14376 21878 14385
rect 21822 14311 21824 14320
rect 21876 14311 21878 14320
rect 21824 14282 21876 14288
rect 21824 12640 21876 12646
rect 21824 12582 21876 12588
rect 21732 12096 21784 12102
rect 21732 12038 21784 12044
rect 21744 11762 21772 12038
rect 21836 11830 21864 12582
rect 21824 11824 21876 11830
rect 21824 11766 21876 11772
rect 21732 11756 21784 11762
rect 21732 11698 21784 11704
rect 21928 11626 21956 17818
rect 22112 17202 22140 19994
rect 22204 19922 22232 20470
rect 22296 20466 22324 21286
rect 22572 21146 22600 21490
rect 22560 21140 22612 21146
rect 22560 21082 22612 21088
rect 22468 21004 22520 21010
rect 22468 20946 22520 20952
rect 22480 20466 22508 20946
rect 22284 20460 22336 20466
rect 22284 20402 22336 20408
rect 22468 20460 22520 20466
rect 22468 20402 22520 20408
rect 22836 20392 22888 20398
rect 22836 20334 22888 20340
rect 22376 20256 22428 20262
rect 22376 20198 22428 20204
rect 22192 19916 22244 19922
rect 22192 19858 22244 19864
rect 22388 19854 22416 20198
rect 22848 19854 22876 20334
rect 22376 19848 22428 19854
rect 22376 19790 22428 19796
rect 22836 19848 22888 19854
rect 22836 19790 22888 19796
rect 22940 19786 22968 29990
rect 23018 29880 23074 29889
rect 23018 29815 23020 29824
rect 23072 29815 23074 29824
rect 23020 29786 23072 29792
rect 23020 29164 23072 29170
rect 23020 29106 23072 29112
rect 23032 28150 23060 29106
rect 23020 28144 23072 28150
rect 23020 28086 23072 28092
rect 23032 27674 23060 28086
rect 23020 27668 23072 27674
rect 23020 27610 23072 27616
rect 23216 27470 23244 30330
rect 23400 29646 23428 31622
rect 23492 30870 23520 31622
rect 23480 30864 23532 30870
rect 23480 30806 23532 30812
rect 23584 30122 23612 32370
rect 23572 30116 23624 30122
rect 23572 30058 23624 30064
rect 23388 29640 23440 29646
rect 23388 29582 23440 29588
rect 23480 29504 23532 29510
rect 23480 29446 23532 29452
rect 23492 28490 23520 29446
rect 23676 28694 23704 32422
rect 23756 32360 23808 32366
rect 23756 32302 23808 32308
rect 23768 31754 23796 32302
rect 23756 31748 23808 31754
rect 23756 31690 23808 31696
rect 23768 29510 23796 31690
rect 23848 31680 23900 31686
rect 23848 31622 23900 31628
rect 23860 30394 23888 31622
rect 24032 31340 24084 31346
rect 24032 31282 24084 31288
rect 23940 31136 23992 31142
rect 23940 31078 23992 31084
rect 23952 30734 23980 31078
rect 23940 30728 23992 30734
rect 23940 30670 23992 30676
rect 23848 30388 23900 30394
rect 23848 30330 23900 30336
rect 24044 29594 24072 31282
rect 24136 30326 24164 32778
rect 24124 30320 24176 30326
rect 24124 30262 24176 30268
rect 24136 30122 24164 30262
rect 24124 30116 24176 30122
rect 24124 30058 24176 30064
rect 24216 29708 24268 29714
rect 24216 29650 24268 29656
rect 23952 29566 24072 29594
rect 24124 29572 24176 29578
rect 23756 29504 23808 29510
rect 23756 29446 23808 29452
rect 23848 29164 23900 29170
rect 23848 29106 23900 29112
rect 23860 28762 23888 29106
rect 23848 28756 23900 28762
rect 23848 28698 23900 28704
rect 23664 28688 23716 28694
rect 23664 28630 23716 28636
rect 23952 28490 23980 29566
rect 24124 29514 24176 29520
rect 24032 29504 24084 29510
rect 24032 29446 24084 29452
rect 23480 28484 23532 28490
rect 23480 28426 23532 28432
rect 23572 28484 23624 28490
rect 23572 28426 23624 28432
rect 23940 28484 23992 28490
rect 23940 28426 23992 28432
rect 23388 28416 23440 28422
rect 23584 28370 23612 28426
rect 23440 28364 23612 28370
rect 23388 28358 23612 28364
rect 23756 28416 23808 28422
rect 23756 28358 23808 28364
rect 23400 28342 23612 28358
rect 23768 28014 23796 28358
rect 23756 28008 23808 28014
rect 23756 27950 23808 27956
rect 23204 27464 23256 27470
rect 23204 27406 23256 27412
rect 23020 27396 23072 27402
rect 23020 27338 23072 27344
rect 23032 26926 23060 27338
rect 23020 26920 23072 26926
rect 23020 26862 23072 26868
rect 23020 26240 23072 26246
rect 23020 26182 23072 26188
rect 23032 25906 23060 26182
rect 23020 25900 23072 25906
rect 23020 25842 23072 25848
rect 23112 25696 23164 25702
rect 23112 25638 23164 25644
rect 23020 24812 23072 24818
rect 23020 24754 23072 24760
rect 23032 24070 23060 24754
rect 23124 24614 23152 25638
rect 23112 24608 23164 24614
rect 23112 24550 23164 24556
rect 23020 24064 23072 24070
rect 23020 24006 23072 24012
rect 23020 23588 23072 23594
rect 23020 23530 23072 23536
rect 23032 20466 23060 23530
rect 23216 22778 23244 27406
rect 23768 27402 23796 27950
rect 23940 27464 23992 27470
rect 23940 27406 23992 27412
rect 23756 27396 23808 27402
rect 23756 27338 23808 27344
rect 23296 27328 23348 27334
rect 23296 27270 23348 27276
rect 23112 22772 23164 22778
rect 23112 22714 23164 22720
rect 23204 22772 23256 22778
rect 23204 22714 23256 22720
rect 23124 22098 23152 22714
rect 23112 22092 23164 22098
rect 23112 22034 23164 22040
rect 23216 21418 23244 22714
rect 23204 21412 23256 21418
rect 23204 21354 23256 21360
rect 23112 21344 23164 21350
rect 23112 21286 23164 21292
rect 23124 20942 23152 21286
rect 23112 20936 23164 20942
rect 23112 20878 23164 20884
rect 23112 20800 23164 20806
rect 23112 20742 23164 20748
rect 23020 20460 23072 20466
rect 23020 20402 23072 20408
rect 22652 19780 22704 19786
rect 22652 19722 22704 19728
rect 22744 19780 22796 19786
rect 22744 19722 22796 19728
rect 22928 19780 22980 19786
rect 22928 19722 22980 19728
rect 22664 19446 22692 19722
rect 22756 19514 22784 19722
rect 23020 19712 23072 19718
rect 23020 19654 23072 19660
rect 22744 19508 22796 19514
rect 22744 19450 22796 19456
rect 22652 19440 22704 19446
rect 22652 19382 22704 19388
rect 22664 17542 22692 19382
rect 22744 18624 22796 18630
rect 22744 18566 22796 18572
rect 22756 18222 22784 18566
rect 22744 18216 22796 18222
rect 22744 18158 22796 18164
rect 22560 17536 22612 17542
rect 22560 17478 22612 17484
rect 22652 17536 22704 17542
rect 22652 17478 22704 17484
rect 22100 17196 22152 17202
rect 22100 17138 22152 17144
rect 22468 16448 22520 16454
rect 22468 16390 22520 16396
rect 22100 15904 22152 15910
rect 22100 15846 22152 15852
rect 22112 12986 22140 15846
rect 22480 15570 22508 16390
rect 22572 16250 22600 17478
rect 22756 17270 22784 18158
rect 22744 17264 22796 17270
rect 22744 17206 22796 17212
rect 22836 16992 22888 16998
rect 22836 16934 22888 16940
rect 22560 16244 22612 16250
rect 22560 16186 22612 16192
rect 22468 15564 22520 15570
rect 22468 15506 22520 15512
rect 22376 15496 22428 15502
rect 22376 15438 22428 15444
rect 22388 14958 22416 15438
rect 22744 15428 22796 15434
rect 22744 15370 22796 15376
rect 22468 15360 22520 15366
rect 22468 15302 22520 15308
rect 22376 14952 22428 14958
rect 22376 14894 22428 14900
rect 22284 14476 22336 14482
rect 22204 14436 22284 14464
rect 22204 14074 22232 14436
rect 22284 14418 22336 14424
rect 22284 14272 22336 14278
rect 22284 14214 22336 14220
rect 22192 14068 22244 14074
rect 22192 14010 22244 14016
rect 22296 13326 22324 14214
rect 22388 14056 22416 14894
rect 22480 14482 22508 15302
rect 22468 14476 22520 14482
rect 22468 14418 22520 14424
rect 22756 14414 22784 15370
rect 22744 14408 22796 14414
rect 22742 14376 22744 14385
rect 22796 14376 22798 14385
rect 22742 14311 22798 14320
rect 22848 14074 22876 16934
rect 23032 16590 23060 19654
rect 23124 18766 23152 20742
rect 23308 20398 23336 27270
rect 23768 26994 23796 27338
rect 23572 26988 23624 26994
rect 23572 26930 23624 26936
rect 23756 26988 23808 26994
rect 23756 26930 23808 26936
rect 23388 26376 23440 26382
rect 23388 26318 23440 26324
rect 23400 25770 23428 26318
rect 23388 25764 23440 25770
rect 23388 25706 23440 25712
rect 23400 25430 23428 25706
rect 23584 25702 23612 26930
rect 23952 25906 23980 27406
rect 23940 25900 23992 25906
rect 23940 25842 23992 25848
rect 23848 25764 23900 25770
rect 23848 25706 23900 25712
rect 23572 25696 23624 25702
rect 23572 25638 23624 25644
rect 23388 25424 23440 25430
rect 23388 25366 23440 25372
rect 23480 25424 23532 25430
rect 23480 25366 23532 25372
rect 23388 25152 23440 25158
rect 23388 25094 23440 25100
rect 23400 23610 23428 25094
rect 23492 24682 23520 25366
rect 23860 25362 23888 25706
rect 23848 25356 23900 25362
rect 23848 25298 23900 25304
rect 23756 25288 23808 25294
rect 23756 25230 23808 25236
rect 23572 25152 23624 25158
rect 23572 25094 23624 25100
rect 23480 24676 23532 24682
rect 23480 24618 23532 24624
rect 23492 24274 23520 24618
rect 23480 24268 23532 24274
rect 23480 24210 23532 24216
rect 23480 24064 23532 24070
rect 23480 24006 23532 24012
rect 23492 23730 23520 24006
rect 23480 23724 23532 23730
rect 23480 23666 23532 23672
rect 23400 23582 23520 23610
rect 23492 23118 23520 23582
rect 23480 23112 23532 23118
rect 23480 23054 23532 23060
rect 23480 22636 23532 22642
rect 23480 22578 23532 22584
rect 23492 22030 23520 22578
rect 23584 22574 23612 25094
rect 23768 24614 23796 25230
rect 23860 24818 23888 25298
rect 23848 24812 23900 24818
rect 23848 24754 23900 24760
rect 23664 24608 23716 24614
rect 23664 24550 23716 24556
rect 23756 24608 23808 24614
rect 23756 24550 23808 24556
rect 23572 22568 23624 22574
rect 23572 22510 23624 22516
rect 23676 22234 23704 24550
rect 23768 23730 23796 24550
rect 23860 23866 23888 24754
rect 23848 23860 23900 23866
rect 23848 23802 23900 23808
rect 23756 23724 23808 23730
rect 23756 23666 23808 23672
rect 23756 23044 23808 23050
rect 23756 22986 23808 22992
rect 23768 22778 23796 22986
rect 23756 22772 23808 22778
rect 23756 22714 23808 22720
rect 23664 22228 23716 22234
rect 23584 22188 23664 22216
rect 23480 22024 23532 22030
rect 23400 21984 23480 22012
rect 23400 21622 23428 21984
rect 23480 21966 23532 21972
rect 23480 21888 23532 21894
rect 23480 21830 23532 21836
rect 23388 21616 23440 21622
rect 23388 21558 23440 21564
rect 23492 20939 23520 21830
rect 23584 21554 23612 22188
rect 23664 22170 23716 22176
rect 23676 22098 23704 22170
rect 23664 22092 23716 22098
rect 23664 22034 23716 22040
rect 23848 22092 23900 22098
rect 23848 22034 23900 22040
rect 23664 21616 23716 21622
rect 23664 21558 23716 21564
rect 23572 21548 23624 21554
rect 23572 21490 23624 21496
rect 23676 21078 23704 21558
rect 23664 21072 23716 21078
rect 23664 21014 23716 21020
rect 23477 20933 23529 20939
rect 23477 20875 23529 20881
rect 23572 20936 23624 20942
rect 23624 20896 23704 20924
rect 23572 20878 23624 20884
rect 23572 20596 23624 20602
rect 23572 20538 23624 20544
rect 23296 20392 23348 20398
rect 23296 20334 23348 20340
rect 23480 20324 23532 20330
rect 23480 20266 23532 20272
rect 23388 19848 23440 19854
rect 23492 19825 23520 20266
rect 23584 19854 23612 20538
rect 23676 20534 23704 20896
rect 23664 20528 23716 20534
rect 23664 20470 23716 20476
rect 23662 20088 23718 20097
rect 23662 20023 23664 20032
rect 23716 20023 23718 20032
rect 23664 19994 23716 20000
rect 23860 19922 23888 22034
rect 24044 21690 24072 29446
rect 24136 29170 24164 29514
rect 24228 29170 24256 29650
rect 24109 29164 24164 29170
rect 24161 29124 24164 29164
rect 24216 29164 24268 29170
rect 24109 29106 24161 29112
rect 24216 29106 24268 29112
rect 24320 28994 24348 36042
rect 24400 35692 24452 35698
rect 24400 35634 24452 35640
rect 24412 35290 24440 35634
rect 24400 35284 24452 35290
rect 24400 35226 24452 35232
rect 24400 35080 24452 35086
rect 24400 35022 24452 35028
rect 24412 33930 24440 35022
rect 24400 33924 24452 33930
rect 24400 33866 24452 33872
rect 24400 33312 24452 33318
rect 24400 33254 24452 33260
rect 24412 32230 24440 33254
rect 24400 32224 24452 32230
rect 24400 32166 24452 32172
rect 24412 31754 24440 32166
rect 24400 31748 24452 31754
rect 24400 31690 24452 31696
rect 24136 28966 24348 28994
rect 24400 29028 24452 29034
rect 24400 28970 24452 28976
rect 24136 26586 24164 28966
rect 24216 28076 24268 28082
rect 24216 28018 24268 28024
rect 24228 27334 24256 28018
rect 24412 27470 24440 28970
rect 24400 27464 24452 27470
rect 24400 27406 24452 27412
rect 24216 27328 24268 27334
rect 24216 27270 24268 27276
rect 24124 26580 24176 26586
rect 24124 26522 24176 26528
rect 24228 26450 24256 27270
rect 24308 26784 24360 26790
rect 24308 26726 24360 26732
rect 24216 26444 24268 26450
rect 24216 26386 24268 26392
rect 24320 26382 24348 26726
rect 24308 26376 24360 26382
rect 24308 26318 24360 26324
rect 24400 26308 24452 26314
rect 24400 26250 24452 26256
rect 24412 25838 24440 26250
rect 24400 25832 24452 25838
rect 24228 25792 24400 25820
rect 24124 25220 24176 25226
rect 24124 25162 24176 25168
rect 24136 24274 24164 25162
rect 24228 24313 24256 25792
rect 24400 25774 24452 25780
rect 24400 25288 24452 25294
rect 24400 25230 24452 25236
rect 24412 24954 24440 25230
rect 24308 24948 24360 24954
rect 24308 24890 24360 24896
rect 24400 24948 24452 24954
rect 24400 24890 24452 24896
rect 24320 24324 24348 24890
rect 24320 24313 24440 24324
rect 24214 24304 24270 24313
rect 24124 24268 24176 24274
rect 24320 24304 24454 24313
rect 24320 24296 24398 24304
rect 24214 24239 24270 24248
rect 24398 24239 24454 24248
rect 24124 24210 24176 24216
rect 24228 24154 24256 24239
rect 24136 24126 24256 24154
rect 24136 22710 24164 24126
rect 24216 24064 24268 24070
rect 24308 24064 24360 24070
rect 24216 24006 24268 24012
rect 24306 24032 24308 24041
rect 24360 24032 24362 24041
rect 24124 22704 24176 22710
rect 24124 22646 24176 22652
rect 24032 21684 24084 21690
rect 24032 21626 24084 21632
rect 24124 21344 24176 21350
rect 24124 21286 24176 21292
rect 24136 21010 24164 21286
rect 24124 21004 24176 21010
rect 24124 20946 24176 20952
rect 24228 20584 24256 24006
rect 24306 23967 24362 23976
rect 24412 23730 24440 24239
rect 24504 24018 24532 37334
rect 25240 36922 25268 37402
rect 25504 37392 25556 37398
rect 25872 37392 25924 37398
rect 25556 37340 25872 37346
rect 25504 37334 25924 37340
rect 25516 37318 25912 37334
rect 25412 37256 25464 37262
rect 25412 37198 25464 37204
rect 25228 36916 25280 36922
rect 25228 36858 25280 36864
rect 24768 36780 24820 36786
rect 24768 36722 24820 36728
rect 24780 36020 24808 36722
rect 24952 36576 25004 36582
rect 24952 36518 25004 36524
rect 24860 36032 24912 36038
rect 24780 35992 24860 36020
rect 24780 35834 24808 35992
rect 24860 35974 24912 35980
rect 24768 35828 24820 35834
rect 24768 35770 24820 35776
rect 24676 34944 24728 34950
rect 24676 34886 24728 34892
rect 24768 34944 24820 34950
rect 24768 34886 24820 34892
rect 24688 34610 24716 34886
rect 24676 34604 24728 34610
rect 24676 34546 24728 34552
rect 24780 34066 24808 34886
rect 24860 34604 24912 34610
rect 24860 34546 24912 34552
rect 24768 34060 24820 34066
rect 24768 34002 24820 34008
rect 24872 33998 24900 34546
rect 24860 33992 24912 33998
rect 24860 33934 24912 33940
rect 24860 33516 24912 33522
rect 24860 33458 24912 33464
rect 24676 33448 24728 33454
rect 24676 33390 24728 33396
rect 24688 33046 24716 33390
rect 24872 33386 24900 33458
rect 24860 33380 24912 33386
rect 24860 33322 24912 33328
rect 24676 33040 24728 33046
rect 24676 32982 24728 32988
rect 24676 32904 24728 32910
rect 24676 32846 24728 32852
rect 24688 32570 24716 32846
rect 24860 32836 24912 32842
rect 24860 32778 24912 32784
rect 24676 32564 24728 32570
rect 24676 32506 24728 32512
rect 24872 32366 24900 32778
rect 24860 32360 24912 32366
rect 24860 32302 24912 32308
rect 24584 31884 24636 31890
rect 24584 31826 24636 31832
rect 24596 31482 24624 31826
rect 24584 31476 24636 31482
rect 24584 31418 24636 31424
rect 24676 31408 24728 31414
rect 24676 31350 24728 31356
rect 24584 30252 24636 30258
rect 24584 30194 24636 30200
rect 24596 29510 24624 30194
rect 24688 29714 24716 31350
rect 24768 30116 24820 30122
rect 24768 30058 24820 30064
rect 24676 29708 24728 29714
rect 24676 29650 24728 29656
rect 24584 29504 24636 29510
rect 24584 29446 24636 29452
rect 24596 29102 24624 29446
rect 24584 29096 24636 29102
rect 24584 29038 24636 29044
rect 24596 28966 24624 29038
rect 24584 28960 24636 28966
rect 24584 28902 24636 28908
rect 24688 27146 24716 29650
rect 24780 29646 24808 30058
rect 24768 29640 24820 29646
rect 24768 29582 24820 29588
rect 24768 29300 24820 29306
rect 24768 29242 24820 29248
rect 24780 28422 24808 29242
rect 24768 28416 24820 28422
rect 24768 28358 24820 28364
rect 24768 28076 24820 28082
rect 24768 28018 24820 28024
rect 24780 27606 24808 28018
rect 24768 27600 24820 27606
rect 24768 27542 24820 27548
rect 24596 27118 24716 27146
rect 24596 26994 24624 27118
rect 24676 27056 24728 27062
rect 24780 27044 24808 27542
rect 24872 27130 24900 32302
rect 24964 31346 24992 36518
rect 25424 36310 25452 37198
rect 25516 36650 25544 37318
rect 25504 36644 25556 36650
rect 25504 36586 25556 36592
rect 25412 36304 25464 36310
rect 25412 36246 25464 36252
rect 25884 36174 25912 37318
rect 27620 37324 27672 37330
rect 27620 37266 27672 37272
rect 26424 37256 26476 37262
rect 26424 37198 26476 37204
rect 26436 37126 26464 37198
rect 26976 37188 27028 37194
rect 26976 37130 27028 37136
rect 26332 37120 26384 37126
rect 26332 37062 26384 37068
rect 26424 37120 26476 37126
rect 26424 37062 26476 37068
rect 26240 36712 26292 36718
rect 26240 36654 26292 36660
rect 26252 36530 26280 36654
rect 26344 36650 26372 37062
rect 26332 36644 26384 36650
rect 26332 36586 26384 36592
rect 26068 36502 26280 36530
rect 26068 36378 26096 36502
rect 26056 36372 26108 36378
rect 26056 36314 26108 36320
rect 26240 36372 26292 36378
rect 26240 36314 26292 36320
rect 25044 36168 25096 36174
rect 25044 36110 25096 36116
rect 25872 36168 25924 36174
rect 25872 36110 25924 36116
rect 25056 33386 25084 36110
rect 26148 35828 26200 35834
rect 26148 35770 26200 35776
rect 25320 35692 25372 35698
rect 25320 35634 25372 35640
rect 25332 35290 25360 35634
rect 25412 35624 25464 35630
rect 25412 35566 25464 35572
rect 25320 35284 25372 35290
rect 25320 35226 25372 35232
rect 25332 34610 25360 35226
rect 25320 34604 25372 34610
rect 25320 34546 25372 34552
rect 25044 33380 25096 33386
rect 25044 33322 25096 33328
rect 25056 32298 25084 33322
rect 25228 32904 25280 32910
rect 25228 32846 25280 32852
rect 25240 32502 25268 32846
rect 25228 32496 25280 32502
rect 25228 32438 25280 32444
rect 25424 32348 25452 35566
rect 26160 35086 26188 35770
rect 25504 35080 25556 35086
rect 25504 35022 25556 35028
rect 25688 35080 25740 35086
rect 25688 35022 25740 35028
rect 26148 35080 26200 35086
rect 26148 35022 26200 35028
rect 25516 34066 25544 35022
rect 25596 34196 25648 34202
rect 25596 34138 25648 34144
rect 25504 34060 25556 34066
rect 25504 34002 25556 34008
rect 25516 33454 25544 34002
rect 25608 33454 25636 34138
rect 25504 33448 25556 33454
rect 25504 33390 25556 33396
rect 25596 33448 25648 33454
rect 25596 33390 25648 33396
rect 25608 33114 25636 33390
rect 25596 33108 25648 33114
rect 25596 33050 25648 33056
rect 25424 32320 25636 32348
rect 25044 32292 25096 32298
rect 25044 32234 25096 32240
rect 25320 32224 25372 32230
rect 25320 32166 25372 32172
rect 25332 32026 25360 32166
rect 25320 32020 25372 32026
rect 25320 31962 25372 31968
rect 25044 31952 25096 31958
rect 25044 31894 25096 31900
rect 25056 31754 25084 31894
rect 25056 31726 25176 31754
rect 24952 31340 25004 31346
rect 24952 31282 25004 31288
rect 24952 30864 25004 30870
rect 24952 30806 25004 30812
rect 24964 30122 24992 30806
rect 25044 30184 25096 30190
rect 25044 30126 25096 30132
rect 24952 30116 25004 30122
rect 24952 30058 25004 30064
rect 24964 28966 24992 30058
rect 25056 29782 25084 30126
rect 25044 29776 25096 29782
rect 25044 29718 25096 29724
rect 25056 29170 25084 29718
rect 25044 29164 25096 29170
rect 25044 29106 25096 29112
rect 24952 28960 25004 28966
rect 24952 28902 25004 28908
rect 24952 28212 25004 28218
rect 24952 28154 25004 28160
rect 25044 28212 25096 28218
rect 25044 28154 25096 28160
rect 24964 27470 24992 28154
rect 25056 28082 25084 28154
rect 25044 28076 25096 28082
rect 25044 28018 25096 28024
rect 24952 27464 25004 27470
rect 24952 27406 25004 27412
rect 24860 27124 24912 27130
rect 24860 27066 24912 27072
rect 24728 27016 24808 27044
rect 24676 26998 24728 27004
rect 24964 26994 24992 27406
rect 24584 26988 24636 26994
rect 24584 26930 24636 26936
rect 24952 26988 25004 26994
rect 24952 26930 25004 26936
rect 24596 26432 24624 26930
rect 24596 26404 24808 26432
rect 24584 25900 24636 25906
rect 24584 25842 24636 25848
rect 24596 24188 24624 25842
rect 24780 25650 24808 26404
rect 24780 25622 24900 25650
rect 24872 25498 24900 25622
rect 24768 25492 24820 25498
rect 24768 25434 24820 25440
rect 24860 25492 24912 25498
rect 24860 25434 24912 25440
rect 24676 25288 24728 25294
rect 24676 25230 24728 25236
rect 24688 24886 24716 25230
rect 24676 24880 24728 24886
rect 24676 24822 24728 24828
rect 24676 24200 24728 24206
rect 24596 24160 24676 24188
rect 24676 24142 24728 24148
rect 24504 23990 24716 24018
rect 24400 23724 24452 23730
rect 24400 23666 24452 23672
rect 24688 23610 24716 23990
rect 24504 23582 24716 23610
rect 24308 22568 24360 22574
rect 24308 22510 24360 22516
rect 24320 21593 24348 22510
rect 24400 22160 24452 22166
rect 24400 22102 24452 22108
rect 24412 21622 24440 22102
rect 24400 21616 24452 21622
rect 24306 21584 24362 21593
rect 24400 21558 24452 21564
rect 24306 21519 24308 21528
rect 24360 21519 24362 21528
rect 24308 21490 24360 21496
rect 24136 20556 24256 20584
rect 23940 20460 23992 20466
rect 23940 20402 23992 20408
rect 23848 19916 23900 19922
rect 23848 19858 23900 19864
rect 23572 19848 23624 19854
rect 23388 19790 23440 19796
rect 23478 19816 23534 19825
rect 23296 19168 23348 19174
rect 23296 19110 23348 19116
rect 23308 18902 23336 19110
rect 23296 18896 23348 18902
rect 23296 18838 23348 18844
rect 23112 18760 23164 18766
rect 23112 18702 23164 18708
rect 23296 18624 23348 18630
rect 23296 18566 23348 18572
rect 23308 17678 23336 18566
rect 23400 17678 23428 19790
rect 23572 19790 23624 19796
rect 23478 19751 23534 19760
rect 23480 19712 23532 19718
rect 23480 19654 23532 19660
rect 23492 18358 23520 19654
rect 23662 19408 23718 19417
rect 23860 19378 23888 19858
rect 23952 19854 23980 20402
rect 23940 19848 23992 19854
rect 23940 19790 23992 19796
rect 23662 19343 23718 19352
rect 23756 19372 23808 19378
rect 23572 19236 23624 19242
rect 23572 19178 23624 19184
rect 23584 18970 23612 19178
rect 23572 18964 23624 18970
rect 23572 18906 23624 18912
rect 23572 18624 23624 18630
rect 23572 18566 23624 18572
rect 23480 18352 23532 18358
rect 23480 18294 23532 18300
rect 23584 18290 23612 18566
rect 23676 18426 23704 19343
rect 23756 19314 23808 19320
rect 23848 19372 23900 19378
rect 23848 19314 23900 19320
rect 23768 18952 23796 19314
rect 23848 18964 23900 18970
rect 23768 18924 23848 18952
rect 23848 18906 23900 18912
rect 24136 18698 24164 20556
rect 24216 20460 24268 20466
rect 24216 20402 24268 20408
rect 24228 20058 24256 20402
rect 24216 20052 24268 20058
rect 24216 19994 24268 20000
rect 24504 19938 24532 23582
rect 24676 23248 24728 23254
rect 24676 23190 24728 23196
rect 24584 22636 24636 22642
rect 24584 22578 24636 22584
rect 24596 22030 24624 22578
rect 24688 22166 24716 23190
rect 24780 22642 24808 25434
rect 24860 24744 24912 24750
rect 24860 24686 24912 24692
rect 24872 23866 24900 24686
rect 24950 24168 25006 24177
rect 24950 24103 25006 24112
rect 24860 23860 24912 23866
rect 24860 23802 24912 23808
rect 24964 23798 24992 24103
rect 24952 23792 25004 23798
rect 24952 23734 25004 23740
rect 24952 23588 25004 23594
rect 24952 23530 25004 23536
rect 24768 22636 24820 22642
rect 24768 22578 24820 22584
rect 24676 22160 24728 22166
rect 24676 22102 24728 22108
rect 24964 22098 24992 23530
rect 25044 23112 25096 23118
rect 25044 23054 25096 23060
rect 25056 22778 25084 23054
rect 25044 22772 25096 22778
rect 25044 22714 25096 22720
rect 24952 22092 25004 22098
rect 24952 22034 25004 22040
rect 24584 22024 24636 22030
rect 24584 21966 24636 21972
rect 24860 22024 24912 22030
rect 24860 21966 24912 21972
rect 24584 21344 24636 21350
rect 24584 21286 24636 21292
rect 24412 19910 24532 19938
rect 24306 18864 24362 18873
rect 24306 18799 24308 18808
rect 24360 18799 24362 18808
rect 24308 18770 24360 18776
rect 24124 18692 24176 18698
rect 24124 18634 24176 18640
rect 23664 18420 23716 18426
rect 23664 18362 23716 18368
rect 23572 18284 23624 18290
rect 23572 18226 23624 18232
rect 23756 17808 23808 17814
rect 23756 17750 23808 17756
rect 23296 17672 23348 17678
rect 23296 17614 23348 17620
rect 23388 17672 23440 17678
rect 23388 17614 23440 17620
rect 23768 17202 23796 17750
rect 23756 17196 23808 17202
rect 23756 17138 23808 17144
rect 23020 16584 23072 16590
rect 23020 16526 23072 16532
rect 23756 16584 23808 16590
rect 23756 16526 23808 16532
rect 23204 16448 23256 16454
rect 23204 16390 23256 16396
rect 23480 16448 23532 16454
rect 23480 16390 23532 16396
rect 23216 16182 23244 16390
rect 23204 16176 23256 16182
rect 23204 16118 23256 16124
rect 23492 16114 23520 16390
rect 23480 16108 23532 16114
rect 23480 16050 23532 16056
rect 22928 16040 22980 16046
rect 22928 15982 22980 15988
rect 22940 15570 22968 15982
rect 23572 15904 23624 15910
rect 23572 15846 23624 15852
rect 22928 15564 22980 15570
rect 22928 15506 22980 15512
rect 23584 15502 23612 15846
rect 23768 15706 23796 16526
rect 24412 16454 24440 19910
rect 24492 19848 24544 19854
rect 24492 19790 24544 19796
rect 24504 19310 24532 19790
rect 24492 19304 24544 19310
rect 24492 19246 24544 19252
rect 24504 18766 24532 19246
rect 24492 18760 24544 18766
rect 24492 18702 24544 18708
rect 24596 17882 24624 21286
rect 24872 20806 24900 21966
rect 24952 21004 25004 21010
rect 24952 20946 25004 20952
rect 24860 20800 24912 20806
rect 24860 20742 24912 20748
rect 24964 20534 24992 20946
rect 24952 20528 25004 20534
rect 24952 20470 25004 20476
rect 25044 20460 25096 20466
rect 25044 20402 25096 20408
rect 24768 20052 24820 20058
rect 24768 19994 24820 20000
rect 24780 19922 24808 19994
rect 24768 19916 24820 19922
rect 24768 19858 24820 19864
rect 25056 19854 25084 20402
rect 24860 19848 24912 19854
rect 24860 19790 24912 19796
rect 25044 19848 25096 19854
rect 25044 19790 25096 19796
rect 24872 18970 24900 19790
rect 24860 18964 24912 18970
rect 24860 18906 24912 18912
rect 24676 18896 24728 18902
rect 24676 18838 24728 18844
rect 24584 17876 24636 17882
rect 24584 17818 24636 17824
rect 24688 17678 24716 18838
rect 25056 18766 25084 19790
rect 25044 18760 25096 18766
rect 25044 18702 25096 18708
rect 25148 18630 25176 31726
rect 25228 30660 25280 30666
rect 25228 30602 25280 30608
rect 25240 30258 25268 30602
rect 25412 30592 25464 30598
rect 25412 30534 25464 30540
rect 25228 30252 25280 30258
rect 25228 30194 25280 30200
rect 25320 30252 25372 30258
rect 25320 30194 25372 30200
rect 25240 29850 25268 30194
rect 25228 29844 25280 29850
rect 25228 29786 25280 29792
rect 25228 29708 25280 29714
rect 25228 29650 25280 29656
rect 25240 29238 25268 29650
rect 25332 29646 25360 30194
rect 25424 29714 25452 30534
rect 25412 29708 25464 29714
rect 25412 29650 25464 29656
rect 25320 29640 25372 29646
rect 25320 29582 25372 29588
rect 25228 29232 25280 29238
rect 25228 29174 25280 29180
rect 25240 28082 25268 29174
rect 25228 28076 25280 28082
rect 25228 28018 25280 28024
rect 25504 27532 25556 27538
rect 25504 27474 25556 27480
rect 25410 27160 25466 27169
rect 25228 27124 25280 27130
rect 25410 27095 25466 27104
rect 25228 27066 25280 27072
rect 25240 25838 25268 27066
rect 25424 27062 25452 27095
rect 25412 27056 25464 27062
rect 25318 27024 25374 27033
rect 25412 26998 25464 27004
rect 25516 26994 25544 27474
rect 25318 26959 25320 26968
rect 25372 26959 25374 26968
rect 25504 26988 25556 26994
rect 25320 26930 25372 26936
rect 25504 26930 25556 26936
rect 25412 26852 25464 26858
rect 25412 26794 25464 26800
rect 25320 26512 25372 26518
rect 25320 26454 25372 26460
rect 25228 25832 25280 25838
rect 25228 25774 25280 25780
rect 25228 24880 25280 24886
rect 25228 24822 25280 24828
rect 25240 24274 25268 24822
rect 25228 24268 25280 24274
rect 25228 24210 25280 24216
rect 25332 23662 25360 26454
rect 25320 23656 25372 23662
rect 25320 23598 25372 23604
rect 25424 23118 25452 26794
rect 25516 26058 25544 26930
rect 25608 26908 25636 32320
rect 25700 32026 25728 35022
rect 26160 34746 26188 35022
rect 26148 34740 26200 34746
rect 26148 34682 26200 34688
rect 25872 34604 25924 34610
rect 25872 34546 25924 34552
rect 25884 33522 25912 34546
rect 25964 33992 26016 33998
rect 25964 33934 26016 33940
rect 25976 33658 26004 33934
rect 25964 33652 26016 33658
rect 25964 33594 26016 33600
rect 25780 33516 25832 33522
rect 25780 33458 25832 33464
rect 25872 33516 25924 33522
rect 25872 33458 25924 33464
rect 26056 33516 26108 33522
rect 26056 33458 26108 33464
rect 25792 32842 25820 33458
rect 25884 32978 25912 33458
rect 25872 32972 25924 32978
rect 25872 32914 25924 32920
rect 25780 32836 25832 32842
rect 25780 32778 25832 32784
rect 25792 32434 25820 32778
rect 26068 32434 26096 33458
rect 25780 32428 25832 32434
rect 25780 32370 25832 32376
rect 26056 32428 26108 32434
rect 26056 32370 26108 32376
rect 25688 32020 25740 32026
rect 25688 31962 25740 31968
rect 25792 31754 25820 32370
rect 26160 31822 26188 34682
rect 26252 33114 26280 36314
rect 26436 36174 26464 37062
rect 26988 36378 27016 37130
rect 27632 36786 27660 37266
rect 28632 37256 28684 37262
rect 28632 37198 28684 37204
rect 30288 37256 30340 37262
rect 30288 37198 30340 37204
rect 28264 37188 28316 37194
rect 28264 37130 28316 37136
rect 28276 36854 28304 37130
rect 28264 36848 28316 36854
rect 28264 36790 28316 36796
rect 28644 36786 28672 37198
rect 29736 37188 29788 37194
rect 29736 37130 29788 37136
rect 28816 37120 28868 37126
rect 28816 37062 28868 37068
rect 28828 36922 28856 37062
rect 28816 36916 28868 36922
rect 28816 36858 28868 36864
rect 29644 36916 29696 36922
rect 29644 36858 29696 36864
rect 27620 36780 27672 36786
rect 27620 36722 27672 36728
rect 28632 36780 28684 36786
rect 28632 36722 28684 36728
rect 27528 36576 27580 36582
rect 27528 36518 27580 36524
rect 27712 36576 27764 36582
rect 27712 36518 27764 36524
rect 28644 36530 28672 36722
rect 28908 36576 28960 36582
rect 27540 36378 27568 36518
rect 26976 36372 27028 36378
rect 26976 36314 27028 36320
rect 27528 36372 27580 36378
rect 27528 36314 27580 36320
rect 26424 36168 26476 36174
rect 26424 36110 26476 36116
rect 26332 35692 26384 35698
rect 26332 35634 26384 35640
rect 26344 35018 26372 35634
rect 26436 35222 26464 36110
rect 26792 35692 26844 35698
rect 26792 35634 26844 35640
rect 26516 35624 26568 35630
rect 26516 35566 26568 35572
rect 26424 35216 26476 35222
rect 26424 35158 26476 35164
rect 26424 35080 26476 35086
rect 26424 35022 26476 35028
rect 26528 35034 26556 35566
rect 26608 35080 26660 35086
rect 26528 35028 26608 35034
rect 26528 35022 26660 35028
rect 26332 35012 26384 35018
rect 26332 34954 26384 34960
rect 26436 34950 26464 35022
rect 26528 35006 26648 35022
rect 26424 34944 26476 34950
rect 26424 34886 26476 34892
rect 26436 34678 26464 34886
rect 26424 34672 26476 34678
rect 26424 34614 26476 34620
rect 26240 33108 26292 33114
rect 26240 33050 26292 33056
rect 26436 32978 26464 34614
rect 26528 34610 26556 35006
rect 26804 34950 26832 35634
rect 27540 35630 27568 36314
rect 27724 35834 27752 36518
rect 28644 36502 28764 36530
rect 28908 36518 28960 36524
rect 28264 36032 28316 36038
rect 28264 35974 28316 35980
rect 28632 36032 28684 36038
rect 28632 35974 28684 35980
rect 27712 35828 27764 35834
rect 27712 35770 27764 35776
rect 27528 35624 27580 35630
rect 27528 35566 27580 35572
rect 28172 35556 28224 35562
rect 28172 35498 28224 35504
rect 27252 35488 27304 35494
rect 27252 35430 27304 35436
rect 26976 35012 27028 35018
rect 26976 34954 27028 34960
rect 26792 34944 26844 34950
rect 26792 34886 26844 34892
rect 26516 34604 26568 34610
rect 26884 34604 26936 34610
rect 26516 34546 26568 34552
rect 26804 34564 26884 34592
rect 26528 33998 26556 34546
rect 26516 33992 26568 33998
rect 26516 33934 26568 33940
rect 26528 33046 26556 33934
rect 26516 33040 26568 33046
rect 26516 32982 26568 32988
rect 26424 32972 26476 32978
rect 26424 32914 26476 32920
rect 26332 32904 26384 32910
rect 26332 32846 26384 32852
rect 26344 32570 26372 32846
rect 26332 32564 26384 32570
rect 26332 32506 26384 32512
rect 26700 32428 26752 32434
rect 26700 32370 26752 32376
rect 26516 32020 26568 32026
rect 26516 31962 26568 31968
rect 26148 31816 26200 31822
rect 26148 31758 26200 31764
rect 25792 31748 26016 31754
rect 25792 31726 25964 31748
rect 25964 31690 26016 31696
rect 25688 31680 25740 31686
rect 25688 31622 25740 31628
rect 25700 29782 25728 31622
rect 25780 31340 25832 31346
rect 25780 31282 25832 31288
rect 25688 29776 25740 29782
rect 25688 29718 25740 29724
rect 25792 27878 25820 31282
rect 25872 28960 25924 28966
rect 25872 28902 25924 28908
rect 25884 28558 25912 28902
rect 25872 28552 25924 28558
rect 25872 28494 25924 28500
rect 25780 27872 25832 27878
rect 25780 27814 25832 27820
rect 25688 27328 25740 27334
rect 25688 27270 25740 27276
rect 25700 27169 25728 27270
rect 25686 27160 25742 27169
rect 25686 27095 25742 27104
rect 25792 26994 25820 27814
rect 25884 27674 25912 28494
rect 25976 28218 26004 31690
rect 26056 31408 26108 31414
rect 26056 31350 26108 31356
rect 25964 28212 26016 28218
rect 25964 28154 26016 28160
rect 25964 27872 26016 27878
rect 25964 27814 26016 27820
rect 25872 27668 25924 27674
rect 25872 27610 25924 27616
rect 25780 26988 25832 26994
rect 25780 26930 25832 26936
rect 25688 26920 25740 26926
rect 25608 26880 25688 26908
rect 25688 26862 25740 26868
rect 25976 26602 26004 27814
rect 26068 27130 26096 31350
rect 26424 31340 26476 31346
rect 26424 31282 26476 31288
rect 26332 31204 26384 31210
rect 26332 31146 26384 31152
rect 26240 30728 26292 30734
rect 26240 30670 26292 30676
rect 26148 30592 26200 30598
rect 26148 30534 26200 30540
rect 26160 30258 26188 30534
rect 26252 30394 26280 30670
rect 26344 30666 26372 31146
rect 26332 30660 26384 30666
rect 26332 30602 26384 30608
rect 26240 30388 26292 30394
rect 26240 30330 26292 30336
rect 26148 30252 26200 30258
rect 26148 30194 26200 30200
rect 26148 29572 26200 29578
rect 26148 29514 26200 29520
rect 26160 29306 26188 29514
rect 26148 29300 26200 29306
rect 26148 29242 26200 29248
rect 26056 27124 26108 27130
rect 26056 27066 26108 27072
rect 25976 26574 26188 26602
rect 25516 26036 25728 26058
rect 25516 26030 25596 26036
rect 25648 26030 25728 26036
rect 25596 25978 25648 25984
rect 25504 25968 25556 25974
rect 25608 25947 25636 25978
rect 25504 25910 25556 25916
rect 25516 24818 25544 25910
rect 25596 25696 25648 25702
rect 25596 25638 25648 25644
rect 25504 24812 25556 24818
rect 25504 24754 25556 24760
rect 25516 24206 25544 24754
rect 25504 24200 25556 24206
rect 25504 24142 25556 24148
rect 25608 23712 25636 25638
rect 25700 24154 25728 26030
rect 25872 26036 25924 26042
rect 25872 25978 25924 25984
rect 25884 25906 25912 25978
rect 25872 25900 25924 25906
rect 26056 25900 26108 25906
rect 25872 25842 25924 25848
rect 25976 25860 26056 25888
rect 25870 25800 25926 25809
rect 25870 25735 25872 25744
rect 25924 25735 25926 25744
rect 25872 25706 25924 25712
rect 25872 25356 25924 25362
rect 25872 25298 25924 25304
rect 25884 25158 25912 25298
rect 25872 25152 25924 25158
rect 25872 25094 25924 25100
rect 25976 24936 26004 25860
rect 26056 25842 26108 25848
rect 26056 25764 26108 25770
rect 26056 25706 26108 25712
rect 25884 24908 26004 24936
rect 25884 24750 25912 24908
rect 26068 24886 26096 25706
rect 26056 24880 26108 24886
rect 26056 24822 26108 24828
rect 25964 24812 26016 24818
rect 25964 24754 26016 24760
rect 25872 24744 25924 24750
rect 25872 24686 25924 24692
rect 25700 24126 25912 24154
rect 25780 24064 25832 24070
rect 25780 24006 25832 24012
rect 25688 23724 25740 23730
rect 25608 23684 25688 23712
rect 25688 23666 25740 23672
rect 25688 23248 25740 23254
rect 25688 23190 25740 23196
rect 25412 23112 25464 23118
rect 25412 23054 25464 23060
rect 25700 22982 25728 23190
rect 25688 22976 25740 22982
rect 25688 22918 25740 22924
rect 25228 22636 25280 22642
rect 25228 22578 25280 22584
rect 25240 21554 25268 22578
rect 25320 22228 25372 22234
rect 25320 22170 25372 22176
rect 25228 21548 25280 21554
rect 25228 21490 25280 21496
rect 25240 21418 25268 21490
rect 25228 21412 25280 21418
rect 25228 21354 25280 21360
rect 25240 21010 25268 21354
rect 25228 21004 25280 21010
rect 25228 20946 25280 20952
rect 25136 18624 25188 18630
rect 25136 18566 25188 18572
rect 24768 18284 24820 18290
rect 24768 18226 24820 18232
rect 24780 17882 24808 18226
rect 25332 18222 25360 22170
rect 25792 22094 25820 24006
rect 25884 23118 25912 24126
rect 25976 24070 26004 24754
rect 26160 24698 26188 26574
rect 26240 25832 26292 25838
rect 26240 25774 26292 25780
rect 26252 24954 26280 25774
rect 26240 24948 26292 24954
rect 26240 24890 26292 24896
rect 26238 24848 26294 24857
rect 26238 24783 26240 24792
rect 26292 24783 26294 24792
rect 26240 24754 26292 24760
rect 26068 24670 26188 24698
rect 25964 24064 26016 24070
rect 25964 24006 26016 24012
rect 25872 23112 25924 23118
rect 25872 23054 25924 23060
rect 25872 22772 25924 22778
rect 25872 22714 25924 22720
rect 25884 22438 25912 22714
rect 25872 22432 25924 22438
rect 25872 22374 25924 22380
rect 25700 22066 25820 22094
rect 25412 22024 25464 22030
rect 25412 21966 25464 21972
rect 25424 21690 25452 21966
rect 25412 21684 25464 21690
rect 25412 21626 25464 21632
rect 25596 20800 25648 20806
rect 25596 20742 25648 20748
rect 25608 20516 25636 20742
rect 25700 20584 25728 22066
rect 25870 21720 25926 21729
rect 25870 21655 25926 21664
rect 25884 21486 25912 21655
rect 25872 21480 25924 21486
rect 25872 21422 25924 21428
rect 25780 20596 25832 20602
rect 25700 20556 25780 20584
rect 25780 20538 25832 20544
rect 25608 20488 25728 20516
rect 25596 20324 25648 20330
rect 25596 20266 25648 20272
rect 25504 20256 25556 20262
rect 25504 20198 25556 20204
rect 25516 19378 25544 20198
rect 25608 19514 25636 20266
rect 25596 19508 25648 19514
rect 25596 19450 25648 19456
rect 25504 19372 25556 19378
rect 25504 19314 25556 19320
rect 25596 19372 25648 19378
rect 25596 19314 25648 19320
rect 25516 18766 25544 19314
rect 25504 18760 25556 18766
rect 25504 18702 25556 18708
rect 25608 18426 25636 19314
rect 25700 19174 25728 20488
rect 25792 19922 25820 20538
rect 25780 19916 25832 19922
rect 25832 19876 25912 19904
rect 25780 19858 25832 19864
rect 25780 19712 25832 19718
rect 25780 19654 25832 19660
rect 25792 19378 25820 19654
rect 25780 19372 25832 19378
rect 25780 19314 25832 19320
rect 25778 19272 25834 19281
rect 25778 19207 25780 19216
rect 25832 19207 25834 19216
rect 25780 19178 25832 19184
rect 25688 19168 25740 19174
rect 25688 19110 25740 19116
rect 25884 18850 25912 19876
rect 25976 19854 26004 24006
rect 26068 22234 26096 24670
rect 26240 24608 26292 24614
rect 26240 24550 26292 24556
rect 26252 24410 26280 24550
rect 26240 24404 26292 24410
rect 26240 24346 26292 24352
rect 26252 23594 26280 24346
rect 26240 23588 26292 23594
rect 26240 23530 26292 23536
rect 26240 23112 26292 23118
rect 26240 23054 26292 23060
rect 26252 22234 26280 23054
rect 26344 22982 26372 30602
rect 26436 26518 26464 31282
rect 26528 30258 26556 31962
rect 26608 31204 26660 31210
rect 26608 31146 26660 31152
rect 26516 30252 26568 30258
rect 26516 30194 26568 30200
rect 26528 29170 26556 30194
rect 26516 29164 26568 29170
rect 26516 29106 26568 29112
rect 26620 29102 26648 31146
rect 26712 30802 26740 32370
rect 26804 31482 26832 34564
rect 26884 34546 26936 34552
rect 26988 33658 27016 34954
rect 26976 33652 27028 33658
rect 26976 33594 27028 33600
rect 27160 32564 27212 32570
rect 27160 32506 27212 32512
rect 27172 32434 27200 32506
rect 27160 32428 27212 32434
rect 27160 32370 27212 32376
rect 26976 32224 27028 32230
rect 26976 32166 27028 32172
rect 26988 32026 27016 32166
rect 26976 32020 27028 32026
rect 26976 31962 27028 31968
rect 26792 31476 26844 31482
rect 26792 31418 26844 31424
rect 26804 31346 26832 31418
rect 27264 31414 27292 35430
rect 27804 35216 27856 35222
rect 27804 35158 27856 35164
rect 27620 35148 27672 35154
rect 27620 35090 27672 35096
rect 27632 34610 27660 35090
rect 27712 34672 27764 34678
rect 27712 34614 27764 34620
rect 27620 34604 27672 34610
rect 27620 34546 27672 34552
rect 27436 33992 27488 33998
rect 27436 33934 27488 33940
rect 27448 33522 27476 33934
rect 27436 33516 27488 33522
rect 27436 33458 27488 33464
rect 27436 32904 27488 32910
rect 27436 32846 27488 32852
rect 27344 32768 27396 32774
rect 27344 32710 27396 32716
rect 27356 32502 27384 32710
rect 27344 32496 27396 32502
rect 27344 32438 27396 32444
rect 27448 32434 27476 32846
rect 27620 32836 27672 32842
rect 27620 32778 27672 32784
rect 27436 32428 27488 32434
rect 27436 32370 27488 32376
rect 27528 31884 27580 31890
rect 27528 31826 27580 31832
rect 27540 31482 27568 31826
rect 27528 31476 27580 31482
rect 27528 31418 27580 31424
rect 27252 31408 27304 31414
rect 27252 31350 27304 31356
rect 26792 31340 26844 31346
rect 26792 31282 26844 31288
rect 27252 31136 27304 31142
rect 27252 31078 27304 31084
rect 26700 30796 26752 30802
rect 26700 30738 26752 30744
rect 27264 30734 27292 31078
rect 27252 30728 27304 30734
rect 27252 30670 27304 30676
rect 27344 30592 27396 30598
rect 27344 30534 27396 30540
rect 27252 29504 27304 29510
rect 27252 29446 27304 29452
rect 27160 29232 27212 29238
rect 27160 29174 27212 29180
rect 26608 29096 26660 29102
rect 26608 29038 26660 29044
rect 26620 28994 26648 29038
rect 26620 28966 26832 28994
rect 26608 27940 26660 27946
rect 26608 27882 26660 27888
rect 26620 27520 26648 27882
rect 26700 27532 26752 27538
rect 26620 27492 26700 27520
rect 26516 27464 26568 27470
rect 26620 27452 26648 27492
rect 26700 27474 26752 27480
rect 26568 27424 26648 27452
rect 26516 27406 26568 27412
rect 26608 27328 26660 27334
rect 26608 27270 26660 27276
rect 26424 26512 26476 26518
rect 26424 26454 26476 26460
rect 26620 26042 26648 27270
rect 26608 26036 26660 26042
rect 26660 25996 26740 26024
rect 26608 25978 26660 25984
rect 26516 25900 26568 25906
rect 26516 25842 26568 25848
rect 26424 25696 26476 25702
rect 26424 25638 26476 25644
rect 26436 24750 26464 25638
rect 26528 25294 26556 25842
rect 26712 25344 26740 25996
rect 26804 25906 26832 28966
rect 27172 28762 27200 29174
rect 27264 29102 27292 29446
rect 27252 29096 27304 29102
rect 27252 29038 27304 29044
rect 27160 28756 27212 28762
rect 27160 28698 27212 28704
rect 27172 28558 27200 28698
rect 26976 28552 27028 28558
rect 26976 28494 27028 28500
rect 27160 28552 27212 28558
rect 27160 28494 27212 28500
rect 26884 27396 26936 27402
rect 26884 27338 26936 27344
rect 26896 26586 26924 27338
rect 26988 26926 27016 28494
rect 27068 28484 27120 28490
rect 27068 28426 27120 28432
rect 26976 26920 27028 26926
rect 26976 26862 27028 26868
rect 27080 26772 27108 28426
rect 27264 28422 27292 29038
rect 27252 28416 27304 28422
rect 27252 28358 27304 28364
rect 26988 26744 27108 26772
rect 26884 26580 26936 26586
rect 26884 26522 26936 26528
rect 26792 25900 26844 25906
rect 26792 25842 26844 25848
rect 26712 25316 26832 25344
rect 26516 25288 26568 25294
rect 26516 25230 26568 25236
rect 26700 25220 26752 25226
rect 26700 25162 26752 25168
rect 26516 25152 26568 25158
rect 26516 25094 26568 25100
rect 26424 24744 26476 24750
rect 26424 24686 26476 24692
rect 26422 24576 26478 24585
rect 26528 24562 26556 25094
rect 26478 24534 26556 24562
rect 26422 24511 26478 24520
rect 26436 24138 26464 24511
rect 26424 24132 26476 24138
rect 26424 24074 26476 24080
rect 26436 23610 26464 24074
rect 26436 23582 26556 23610
rect 26424 23520 26476 23526
rect 26424 23462 26476 23468
rect 26332 22976 26384 22982
rect 26332 22918 26384 22924
rect 26056 22228 26108 22234
rect 26056 22170 26108 22176
rect 26240 22228 26292 22234
rect 26240 22170 26292 22176
rect 26148 21888 26200 21894
rect 26148 21830 26200 21836
rect 26056 21548 26108 21554
rect 26056 21490 26108 21496
rect 26068 21350 26096 21490
rect 26056 21344 26108 21350
rect 26056 21286 26108 21292
rect 26056 20256 26108 20262
rect 26056 20198 26108 20204
rect 26068 20097 26096 20198
rect 26054 20088 26110 20097
rect 26054 20023 26110 20032
rect 26160 19990 26188 21830
rect 26436 21622 26464 23462
rect 26528 22166 26556 23582
rect 26608 23316 26660 23322
rect 26608 23258 26660 23264
rect 26620 23186 26648 23258
rect 26608 23180 26660 23186
rect 26608 23122 26660 23128
rect 26516 22160 26568 22166
rect 26516 22102 26568 22108
rect 26424 21616 26476 21622
rect 26424 21558 26476 21564
rect 26332 21548 26384 21554
rect 26332 21490 26384 21496
rect 26344 21418 26372 21490
rect 26332 21412 26384 21418
rect 26332 21354 26384 21360
rect 26240 21344 26292 21350
rect 26240 21286 26292 21292
rect 26148 19984 26200 19990
rect 26148 19926 26200 19932
rect 25964 19848 26016 19854
rect 25964 19790 26016 19796
rect 25792 18822 25912 18850
rect 25596 18420 25648 18426
rect 25596 18362 25648 18368
rect 25792 18290 25820 18822
rect 25872 18760 25924 18766
rect 25872 18702 25924 18708
rect 25884 18426 25912 18702
rect 25872 18420 25924 18426
rect 25872 18362 25924 18368
rect 25976 18358 26004 19790
rect 26252 19514 26280 21286
rect 26344 21010 26372 21354
rect 26332 21004 26384 21010
rect 26332 20946 26384 20952
rect 26424 20800 26476 20806
rect 26424 20742 26476 20748
rect 26332 20324 26384 20330
rect 26332 20266 26384 20272
rect 26344 19854 26372 20266
rect 26332 19848 26384 19854
rect 26332 19790 26384 19796
rect 26240 19508 26292 19514
rect 26240 19450 26292 19456
rect 26252 19378 26280 19450
rect 26240 19372 26292 19378
rect 26240 19314 26292 19320
rect 26056 19304 26108 19310
rect 26056 19246 26108 19252
rect 26068 19174 26096 19246
rect 26056 19168 26108 19174
rect 26056 19110 26108 19116
rect 26240 19168 26292 19174
rect 26240 19110 26292 19116
rect 25964 18352 26016 18358
rect 25964 18294 26016 18300
rect 25780 18284 25832 18290
rect 25780 18226 25832 18232
rect 25320 18216 25372 18222
rect 25320 18158 25372 18164
rect 26068 18154 26096 19110
rect 26252 18698 26280 19110
rect 26344 18766 26372 19790
rect 26332 18760 26384 18766
rect 26332 18702 26384 18708
rect 26240 18692 26292 18698
rect 26240 18634 26292 18640
rect 26148 18624 26200 18630
rect 26148 18566 26200 18572
rect 26160 18290 26188 18566
rect 26148 18284 26200 18290
rect 26148 18226 26200 18232
rect 26056 18148 26108 18154
rect 26056 18090 26108 18096
rect 25228 18080 25280 18086
rect 25228 18022 25280 18028
rect 24768 17876 24820 17882
rect 24768 17818 24820 17824
rect 24676 17672 24728 17678
rect 24676 17614 24728 17620
rect 25240 17202 25268 18022
rect 25504 17672 25556 17678
rect 25504 17614 25556 17620
rect 25228 17196 25280 17202
rect 25228 17138 25280 17144
rect 25412 16584 25464 16590
rect 25412 16526 25464 16532
rect 24400 16448 24452 16454
rect 24400 16390 24452 16396
rect 25424 16250 25452 16526
rect 25044 16244 25096 16250
rect 25044 16186 25096 16192
rect 25412 16244 25464 16250
rect 25412 16186 25464 16192
rect 25056 15706 25084 16186
rect 25516 16114 25544 17614
rect 26436 17610 26464 20742
rect 26516 20528 26568 20534
rect 26516 20470 26568 20476
rect 26528 19718 26556 20470
rect 26712 20466 26740 25162
rect 26804 24818 26832 25316
rect 26884 25288 26936 25294
rect 26884 25230 26936 25236
rect 26792 24812 26844 24818
rect 26792 24754 26844 24760
rect 26792 24608 26844 24614
rect 26792 24550 26844 24556
rect 26804 24206 26832 24550
rect 26896 24410 26924 25230
rect 26884 24404 26936 24410
rect 26884 24346 26936 24352
rect 26792 24200 26844 24206
rect 26792 24142 26844 24148
rect 26792 23724 26844 23730
rect 26792 23666 26844 23672
rect 26804 23322 26832 23666
rect 26988 23594 27016 26744
rect 27066 26480 27122 26489
rect 27066 26415 27122 26424
rect 27080 26382 27108 26415
rect 27068 26376 27120 26382
rect 27068 26318 27120 26324
rect 27264 26246 27292 28358
rect 27252 26240 27304 26246
rect 27252 26182 27304 26188
rect 27068 25288 27120 25294
rect 27068 25230 27120 25236
rect 27080 24614 27108 25230
rect 27252 24744 27304 24750
rect 27252 24686 27304 24692
rect 27068 24608 27120 24614
rect 27068 24550 27120 24556
rect 27264 24274 27292 24686
rect 27252 24268 27304 24274
rect 27252 24210 27304 24216
rect 27160 24200 27212 24206
rect 27160 24142 27212 24148
rect 26976 23588 27028 23594
rect 26976 23530 27028 23536
rect 27172 23526 27200 24142
rect 27252 23724 27304 23730
rect 27252 23666 27304 23672
rect 27160 23520 27212 23526
rect 27160 23462 27212 23468
rect 26792 23316 26844 23322
rect 26792 23258 26844 23264
rect 26804 22438 26832 23258
rect 26884 23112 26936 23118
rect 26884 23054 26936 23060
rect 26896 22574 26924 23054
rect 27068 23044 27120 23050
rect 27068 22986 27120 22992
rect 27080 22642 27108 22986
rect 26976 22636 27028 22642
rect 26976 22578 27028 22584
rect 27068 22636 27120 22642
rect 27068 22578 27120 22584
rect 26884 22568 26936 22574
rect 26884 22510 26936 22516
rect 26792 22432 26844 22438
rect 26792 22374 26844 22380
rect 26804 20942 26832 22374
rect 26988 22216 27016 22578
rect 26988 22188 27108 22216
rect 26884 22160 26936 22166
rect 26936 22108 27016 22114
rect 26884 22102 27016 22108
rect 26896 22086 27016 22102
rect 27080 22098 27108 22188
rect 26792 20936 26844 20942
rect 26792 20878 26844 20884
rect 26804 20534 26832 20878
rect 26792 20528 26844 20534
rect 26792 20470 26844 20476
rect 26700 20460 26752 20466
rect 26700 20402 26752 20408
rect 26884 20460 26936 20466
rect 26884 20402 26936 20408
rect 26896 19990 26924 20402
rect 26884 19984 26936 19990
rect 26884 19926 26936 19932
rect 26516 19712 26568 19718
rect 26516 19654 26568 19660
rect 26988 18766 27016 22086
rect 27068 22092 27120 22098
rect 27172 22094 27200 23462
rect 27264 22982 27292 23666
rect 27252 22976 27304 22982
rect 27252 22918 27304 22924
rect 27356 22710 27384 30534
rect 27632 30410 27660 32778
rect 27724 32756 27752 34614
rect 27816 33998 27844 35158
rect 27896 35080 27948 35086
rect 27896 35022 27948 35028
rect 28080 35080 28132 35086
rect 28080 35022 28132 35028
rect 27908 34746 27936 35022
rect 27988 34944 28040 34950
rect 27988 34886 28040 34892
rect 27896 34740 27948 34746
rect 27896 34682 27948 34688
rect 28000 34678 28028 34886
rect 27988 34672 28040 34678
rect 27988 34614 28040 34620
rect 28092 34406 28120 35022
rect 28184 34950 28212 35498
rect 28172 34944 28224 34950
rect 28172 34886 28224 34892
rect 28184 34610 28212 34886
rect 28172 34604 28224 34610
rect 28172 34546 28224 34552
rect 28080 34400 28132 34406
rect 28080 34342 28132 34348
rect 27804 33992 27856 33998
rect 27804 33934 27856 33940
rect 28172 32768 28224 32774
rect 27724 32728 27844 32756
rect 27540 30382 27660 30410
rect 27540 30190 27568 30382
rect 27816 30258 27844 32728
rect 28172 32710 28224 32716
rect 28184 32434 28212 32710
rect 28172 32428 28224 32434
rect 28172 32370 28224 32376
rect 28184 31822 28212 32370
rect 28172 31816 28224 31822
rect 28172 31758 28224 31764
rect 28276 31210 28304 35974
rect 28540 35828 28592 35834
rect 28540 35770 28592 35776
rect 28448 35692 28500 35698
rect 28448 35634 28500 35640
rect 28356 35624 28408 35630
rect 28356 35566 28408 35572
rect 28264 31204 28316 31210
rect 28264 31146 28316 31152
rect 28080 31136 28132 31142
rect 28080 31078 28132 31084
rect 28092 30802 28120 31078
rect 28368 30802 28396 35566
rect 28460 35494 28488 35634
rect 28448 35488 28500 35494
rect 28448 35430 28500 35436
rect 28460 35018 28488 35430
rect 28552 35086 28580 35770
rect 28644 35290 28672 35974
rect 28736 35766 28764 36502
rect 28816 36372 28868 36378
rect 28816 36314 28868 36320
rect 28828 36242 28856 36314
rect 28920 36310 28948 36518
rect 28908 36304 28960 36310
rect 28908 36246 28960 36252
rect 28816 36236 28868 36242
rect 28816 36178 28868 36184
rect 28724 35760 28776 35766
rect 28724 35702 28776 35708
rect 28632 35284 28684 35290
rect 28632 35226 28684 35232
rect 28828 35154 28856 36178
rect 29656 36174 29684 36858
rect 29748 36786 29776 37130
rect 29736 36780 29788 36786
rect 29736 36722 29788 36728
rect 29828 36780 29880 36786
rect 29828 36722 29880 36728
rect 29644 36168 29696 36174
rect 29644 36110 29696 36116
rect 29748 35834 29776 36722
rect 29736 35828 29788 35834
rect 29736 35770 29788 35776
rect 29840 35290 29868 36722
rect 30196 36712 30248 36718
rect 30196 36654 30248 36660
rect 30208 36174 30236 36654
rect 30300 36310 30328 37198
rect 30472 37120 30524 37126
rect 34440 37108 34468 39222
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 35808 37256 35860 37262
rect 35808 37198 35860 37204
rect 34520 37120 34572 37126
rect 34440 37080 34520 37108
rect 30472 37062 30524 37068
rect 34520 37062 34572 37068
rect 30484 36786 30512 37062
rect 30472 36780 30524 36786
rect 30472 36722 30524 36728
rect 30932 36712 30984 36718
rect 30932 36654 30984 36660
rect 30380 36644 30432 36650
rect 30380 36586 30432 36592
rect 30288 36304 30340 36310
rect 30288 36246 30340 36252
rect 30196 36168 30248 36174
rect 30196 36110 30248 36116
rect 30288 36032 30340 36038
rect 30288 35974 30340 35980
rect 30300 35834 30328 35974
rect 30288 35828 30340 35834
rect 30288 35770 30340 35776
rect 30392 35698 30420 36586
rect 30944 36378 30972 36654
rect 32496 36644 32548 36650
rect 32496 36586 32548 36592
rect 30932 36372 30984 36378
rect 30932 36314 30984 36320
rect 31576 36372 31628 36378
rect 31576 36314 31628 36320
rect 31208 36168 31260 36174
rect 31208 36110 31260 36116
rect 30380 35692 30432 35698
rect 30380 35634 30432 35640
rect 29828 35284 29880 35290
rect 29828 35226 29880 35232
rect 28816 35148 28868 35154
rect 28816 35090 28868 35096
rect 30932 35148 30984 35154
rect 30932 35090 30984 35096
rect 28540 35080 28592 35086
rect 28540 35022 28592 35028
rect 30288 35080 30340 35086
rect 30288 35022 30340 35028
rect 30380 35080 30432 35086
rect 30380 35022 30432 35028
rect 28448 35012 28500 35018
rect 28448 34954 28500 34960
rect 28552 34762 28580 35022
rect 29736 34944 29788 34950
rect 29736 34886 29788 34892
rect 30196 34944 30248 34950
rect 30196 34886 30248 34892
rect 28460 34734 28580 34762
rect 28460 34202 28488 34734
rect 28540 34672 28592 34678
rect 28540 34614 28592 34620
rect 28448 34196 28500 34202
rect 28448 34138 28500 34144
rect 28448 33516 28500 33522
rect 28448 33458 28500 33464
rect 28460 32842 28488 33458
rect 28552 33114 28580 34614
rect 29276 34604 29328 34610
rect 29276 34546 29328 34552
rect 29460 34604 29512 34610
rect 29460 34546 29512 34552
rect 28632 34400 28684 34406
rect 28632 34342 28684 34348
rect 28816 34400 28868 34406
rect 28816 34342 28868 34348
rect 28644 33522 28672 34342
rect 28828 34066 28856 34342
rect 28816 34060 28868 34066
rect 28816 34002 28868 34008
rect 28724 33924 28776 33930
rect 28724 33866 28776 33872
rect 28632 33516 28684 33522
rect 28632 33458 28684 33464
rect 28736 33386 28764 33866
rect 29288 33590 29316 34546
rect 29276 33584 29328 33590
rect 29276 33526 29328 33532
rect 29472 33522 29500 34546
rect 29644 34196 29696 34202
rect 29644 34138 29696 34144
rect 29656 34066 29684 34138
rect 29644 34060 29696 34066
rect 29644 34002 29696 34008
rect 29092 33516 29144 33522
rect 29092 33458 29144 33464
rect 29460 33516 29512 33522
rect 29460 33458 29512 33464
rect 29000 33448 29052 33454
rect 29000 33390 29052 33396
rect 28724 33380 28776 33386
rect 28724 33322 28776 33328
rect 28540 33108 28592 33114
rect 28540 33050 28592 33056
rect 29012 32910 29040 33390
rect 29104 32978 29132 33458
rect 29656 32978 29684 34002
rect 29092 32972 29144 32978
rect 29092 32914 29144 32920
rect 29644 32972 29696 32978
rect 29644 32914 29696 32920
rect 29000 32904 29052 32910
rect 29000 32846 29052 32852
rect 28448 32836 28500 32842
rect 28448 32778 28500 32784
rect 28540 32768 28592 32774
rect 28540 32710 28592 32716
rect 28552 32570 28580 32710
rect 29012 32570 29040 32846
rect 28540 32564 28592 32570
rect 28540 32506 28592 32512
rect 29000 32564 29052 32570
rect 29000 32506 29052 32512
rect 28448 32292 28500 32298
rect 28448 32234 28500 32240
rect 28460 31822 28488 32234
rect 28908 32224 28960 32230
rect 28908 32166 28960 32172
rect 28448 31816 28500 31822
rect 28448 31758 28500 31764
rect 28540 31748 28592 31754
rect 28540 31690 28592 31696
rect 28552 31346 28580 31690
rect 28724 31680 28776 31686
rect 28724 31622 28776 31628
rect 28540 31340 28592 31346
rect 28540 31282 28592 31288
rect 28080 30796 28132 30802
rect 28080 30738 28132 30744
rect 28356 30796 28408 30802
rect 28356 30738 28408 30744
rect 28080 30320 28132 30326
rect 28080 30262 28132 30268
rect 27804 30252 27856 30258
rect 27620 30218 27672 30224
rect 27528 30184 27580 30190
rect 27804 30194 27856 30200
rect 27620 30160 27672 30166
rect 27528 30126 27580 30132
rect 27632 29306 27660 30160
rect 27620 29300 27672 29306
rect 27620 29242 27672 29248
rect 27632 28762 27660 29242
rect 27712 29028 27764 29034
rect 27712 28970 27764 28976
rect 27620 28756 27672 28762
rect 27620 28698 27672 28704
rect 27528 28688 27580 28694
rect 27528 28630 27580 28636
rect 27436 27872 27488 27878
rect 27434 27840 27436 27849
rect 27488 27840 27490 27849
rect 27434 27775 27490 27784
rect 27436 27464 27488 27470
rect 27436 27406 27488 27412
rect 27448 27033 27476 27406
rect 27434 27024 27490 27033
rect 27540 26994 27568 28630
rect 27724 28082 27752 28970
rect 27816 28626 27844 30194
rect 28092 30054 28120 30262
rect 28172 30184 28224 30190
rect 28172 30126 28224 30132
rect 28264 30184 28316 30190
rect 28264 30126 28316 30132
rect 28080 30048 28132 30054
rect 28080 29990 28132 29996
rect 28080 29640 28132 29646
rect 28080 29582 28132 29588
rect 28092 29306 28120 29582
rect 28184 29510 28212 30126
rect 28276 29889 28304 30126
rect 28262 29880 28318 29889
rect 28262 29815 28318 29824
rect 28172 29504 28224 29510
rect 28172 29446 28224 29452
rect 28080 29300 28132 29306
rect 28080 29242 28132 29248
rect 28368 28994 28396 30738
rect 28552 30734 28580 31282
rect 28540 30728 28592 30734
rect 28540 30670 28592 30676
rect 28540 30388 28592 30394
rect 28540 30330 28592 30336
rect 28448 30252 28500 30258
rect 28448 30194 28500 30200
rect 28460 29034 28488 30194
rect 28552 29238 28580 30330
rect 28632 30048 28684 30054
rect 28632 29990 28684 29996
rect 28540 29232 28592 29238
rect 28540 29174 28592 29180
rect 28276 28966 28396 28994
rect 28448 29028 28500 29034
rect 28448 28970 28500 28976
rect 27804 28620 27856 28626
rect 27804 28562 27856 28568
rect 28172 28552 28224 28558
rect 28078 28520 28134 28529
rect 28172 28494 28224 28500
rect 28078 28455 28134 28464
rect 27988 28416 28040 28422
rect 27988 28358 28040 28364
rect 27712 28076 27764 28082
rect 27712 28018 27764 28024
rect 27620 27940 27672 27946
rect 27620 27882 27672 27888
rect 27434 26959 27490 26968
rect 27528 26988 27580 26994
rect 27528 26930 27580 26936
rect 27436 26920 27488 26926
rect 27436 26862 27488 26868
rect 27448 25974 27476 26862
rect 27528 26784 27580 26790
rect 27528 26726 27580 26732
rect 27540 26382 27568 26726
rect 27528 26376 27580 26382
rect 27528 26318 27580 26324
rect 27436 25968 27488 25974
rect 27436 25910 27488 25916
rect 27632 25362 27660 27882
rect 27894 27704 27950 27713
rect 27894 27639 27896 27648
rect 27948 27639 27950 27648
rect 27896 27610 27948 27616
rect 28000 27402 28028 28358
rect 28092 28014 28120 28455
rect 28184 28218 28212 28494
rect 28172 28212 28224 28218
rect 28172 28154 28224 28160
rect 28172 28076 28224 28082
rect 28172 28018 28224 28024
rect 28080 28008 28132 28014
rect 28080 27950 28132 27956
rect 28184 27606 28212 28018
rect 28080 27600 28132 27606
rect 28078 27568 28080 27577
rect 28172 27600 28224 27606
rect 28132 27568 28134 27577
rect 28172 27542 28224 27548
rect 28078 27503 28134 27512
rect 27712 27396 27764 27402
rect 27712 27338 27764 27344
rect 27988 27396 28040 27402
rect 27988 27338 28040 27344
rect 27724 26586 27752 27338
rect 27712 26580 27764 26586
rect 27712 26522 27764 26528
rect 27804 26580 27856 26586
rect 27804 26522 27856 26528
rect 27816 26382 27844 26522
rect 27804 26376 27856 26382
rect 27804 26318 27856 26324
rect 27816 25770 27844 26318
rect 28000 25974 28028 27338
rect 28080 26988 28132 26994
rect 28080 26930 28132 26936
rect 28092 26897 28120 26930
rect 28078 26888 28134 26897
rect 28078 26823 28134 26832
rect 28172 26512 28224 26518
rect 28172 26454 28224 26460
rect 27988 25968 28040 25974
rect 27988 25910 28040 25916
rect 27804 25764 27856 25770
rect 27804 25706 27856 25712
rect 27620 25356 27672 25362
rect 27620 25298 27672 25304
rect 28080 25288 28132 25294
rect 28080 25230 28132 25236
rect 27620 25152 27672 25158
rect 27620 25094 27672 25100
rect 27528 24880 27580 24886
rect 27528 24822 27580 24828
rect 27436 24336 27488 24342
rect 27436 24278 27488 24284
rect 27448 24018 27476 24278
rect 27540 24206 27568 24822
rect 27528 24200 27580 24206
rect 27528 24142 27580 24148
rect 27632 24018 27660 25094
rect 28092 24818 28120 25230
rect 28080 24812 28132 24818
rect 28080 24754 28132 24760
rect 27988 24336 28040 24342
rect 27986 24304 27988 24313
rect 28040 24304 28042 24313
rect 27986 24239 28042 24248
rect 27448 23990 27660 24018
rect 27448 23730 27476 23990
rect 28184 23905 28212 26454
rect 28276 25809 28304 28966
rect 28446 28928 28502 28937
rect 28446 28863 28502 28872
rect 28460 27962 28488 28863
rect 28552 28490 28580 29174
rect 28540 28484 28592 28490
rect 28540 28426 28592 28432
rect 28460 27934 28580 27962
rect 28448 27872 28500 27878
rect 28446 27840 28448 27849
rect 28500 27840 28502 27849
rect 28446 27775 28502 27784
rect 28446 27704 28502 27713
rect 28446 27639 28448 27648
rect 28500 27639 28502 27648
rect 28448 27610 28500 27616
rect 28552 27606 28580 27934
rect 28540 27600 28592 27606
rect 28540 27542 28592 27548
rect 28356 27328 28408 27334
rect 28356 27270 28408 27276
rect 28540 27328 28592 27334
rect 28540 27270 28592 27276
rect 28368 26926 28396 27270
rect 28448 27056 28500 27062
rect 28448 26998 28500 27004
rect 28356 26920 28408 26926
rect 28356 26862 28408 26868
rect 28368 26194 28396 26862
rect 28460 26790 28488 26998
rect 28448 26784 28500 26790
rect 28448 26726 28500 26732
rect 28552 26382 28580 27270
rect 28540 26376 28592 26382
rect 28540 26318 28592 26324
rect 28368 26166 28488 26194
rect 28356 26036 28408 26042
rect 28356 25978 28408 25984
rect 28262 25800 28318 25809
rect 28262 25735 28318 25744
rect 28276 24886 28304 25735
rect 28264 24880 28316 24886
rect 28264 24822 28316 24828
rect 28170 23896 28226 23905
rect 28080 23860 28132 23866
rect 28170 23831 28226 23840
rect 28080 23802 28132 23808
rect 27436 23724 27488 23730
rect 27436 23666 27488 23672
rect 27436 23588 27488 23594
rect 27436 23530 27488 23536
rect 27344 22704 27396 22710
rect 27344 22646 27396 22652
rect 27344 22568 27396 22574
rect 27344 22510 27396 22516
rect 27172 22066 27292 22094
rect 27068 22034 27120 22040
rect 27080 21622 27108 22034
rect 27160 21888 27212 21894
rect 27160 21830 27212 21836
rect 27068 21616 27120 21622
rect 27068 21558 27120 21564
rect 27068 21004 27120 21010
rect 27068 20946 27120 20952
rect 27080 20466 27108 20946
rect 27068 20460 27120 20466
rect 27068 20402 27120 20408
rect 26792 18760 26844 18766
rect 26792 18702 26844 18708
rect 26976 18760 27028 18766
rect 26976 18702 27028 18708
rect 26804 18358 26832 18702
rect 26976 18624 27028 18630
rect 26976 18566 27028 18572
rect 26988 18426 27016 18566
rect 26976 18420 27028 18426
rect 26976 18362 27028 18368
rect 26792 18352 26844 18358
rect 26792 18294 26844 18300
rect 26804 17814 26832 18294
rect 26792 17808 26844 17814
rect 26792 17750 26844 17756
rect 27172 17678 27200 21830
rect 27264 17746 27292 22066
rect 27356 21554 27384 22510
rect 27344 21548 27396 21554
rect 27344 21490 27396 21496
rect 27448 20641 27476 23530
rect 27988 23520 28040 23526
rect 27988 23462 28040 23468
rect 27804 23316 27856 23322
rect 27804 23258 27856 23264
rect 27528 23180 27580 23186
rect 27528 23122 27580 23128
rect 27540 22642 27568 23122
rect 27816 23118 27844 23258
rect 28000 23118 28028 23462
rect 28092 23254 28120 23802
rect 28080 23248 28132 23254
rect 28080 23190 28132 23196
rect 28368 23186 28396 25978
rect 28356 23180 28408 23186
rect 28356 23122 28408 23128
rect 27804 23112 27856 23118
rect 27724 23072 27804 23100
rect 27528 22636 27580 22642
rect 27528 22578 27580 22584
rect 27528 22432 27580 22438
rect 27528 22374 27580 22380
rect 27540 22098 27568 22374
rect 27724 22166 27752 23072
rect 27804 23054 27856 23060
rect 27988 23112 28040 23118
rect 27988 23054 28040 23060
rect 27804 22432 27856 22438
rect 27804 22374 27856 22380
rect 28264 22432 28316 22438
rect 28264 22374 28316 22380
rect 27712 22160 27764 22166
rect 27712 22102 27764 22108
rect 27528 22092 27580 22098
rect 27528 22034 27580 22040
rect 27620 21140 27672 21146
rect 27620 21082 27672 21088
rect 27712 21140 27764 21146
rect 27712 21082 27764 21088
rect 27434 20632 27490 20641
rect 27434 20567 27490 20576
rect 27632 20244 27660 21082
rect 27724 20534 27752 21082
rect 27712 20528 27764 20534
rect 27712 20470 27764 20476
rect 27712 20256 27764 20262
rect 27632 20216 27712 20244
rect 27712 20198 27764 20204
rect 27342 19680 27398 19689
rect 27342 19615 27398 19624
rect 27356 19446 27384 19615
rect 27344 19440 27396 19446
rect 27344 19382 27396 19388
rect 27252 17740 27304 17746
rect 27252 17682 27304 17688
rect 27160 17672 27212 17678
rect 27160 17614 27212 17620
rect 26424 17604 26476 17610
rect 26424 17546 26476 17552
rect 27816 17542 27844 22374
rect 28172 22228 28224 22234
rect 28172 22170 28224 22176
rect 27988 22024 28040 22030
rect 27988 21966 28040 21972
rect 27896 21888 27948 21894
rect 27896 21830 27948 21836
rect 27908 21690 27936 21830
rect 28000 21690 28028 21966
rect 27896 21684 27948 21690
rect 27896 21626 27948 21632
rect 27988 21684 28040 21690
rect 27988 21626 28040 21632
rect 27896 21344 27948 21350
rect 27896 21286 27948 21292
rect 27908 21010 27936 21286
rect 27896 21004 27948 21010
rect 27896 20946 27948 20952
rect 27896 20868 27948 20874
rect 27896 20810 27948 20816
rect 28080 20868 28132 20874
rect 28080 20810 28132 20816
rect 27908 19242 27936 20810
rect 27986 20632 28042 20641
rect 27986 20567 28042 20576
rect 28000 20534 28028 20567
rect 27988 20528 28040 20534
rect 27988 20470 28040 20476
rect 28092 20398 28120 20810
rect 28080 20392 28132 20398
rect 28080 20334 28132 20340
rect 27986 19816 28042 19825
rect 27986 19751 28042 19760
rect 27896 19236 27948 19242
rect 27896 19178 27948 19184
rect 27908 18970 27936 19178
rect 27896 18964 27948 18970
rect 27896 18906 27948 18912
rect 28000 18086 28028 19751
rect 28184 19718 28212 22170
rect 28276 22098 28304 22374
rect 28460 22234 28488 26166
rect 28644 25838 28672 29990
rect 28736 29306 28764 31622
rect 28920 30870 28948 32166
rect 29104 31958 29132 32914
rect 29552 32428 29604 32434
rect 29552 32370 29604 32376
rect 29092 31952 29144 31958
rect 29092 31894 29144 31900
rect 29564 31890 29592 32370
rect 29552 31884 29604 31890
rect 29472 31844 29552 31872
rect 29092 31340 29144 31346
rect 29092 31282 29144 31288
rect 28908 30864 28960 30870
rect 28908 30806 28960 30812
rect 29000 30728 29052 30734
rect 29000 30670 29052 30676
rect 28816 30592 28868 30598
rect 28816 30534 28868 30540
rect 28724 29300 28776 29306
rect 28724 29242 28776 29248
rect 28724 28620 28776 28626
rect 28724 28562 28776 28568
rect 28736 28150 28764 28562
rect 28828 28150 28856 30534
rect 29012 29850 29040 30670
rect 29104 30326 29132 31282
rect 29472 30598 29500 31844
rect 29552 31826 29604 31832
rect 29552 31272 29604 31278
rect 29552 31214 29604 31220
rect 29460 30592 29512 30598
rect 29460 30534 29512 30540
rect 29092 30320 29144 30326
rect 29092 30262 29144 30268
rect 29000 29844 29052 29850
rect 29000 29786 29052 29792
rect 29368 29844 29420 29850
rect 29368 29786 29420 29792
rect 28908 29708 28960 29714
rect 28908 29650 28960 29656
rect 29092 29708 29144 29714
rect 29092 29650 29144 29656
rect 28920 29238 28948 29650
rect 29104 29458 29132 29650
rect 29184 29572 29236 29578
rect 29184 29514 29236 29520
rect 29012 29430 29132 29458
rect 28908 29232 28960 29238
rect 28908 29174 28960 29180
rect 29012 29084 29040 29430
rect 29092 29232 29144 29238
rect 29090 29200 29092 29209
rect 29144 29200 29146 29209
rect 29090 29135 29146 29144
rect 28920 29056 29040 29084
rect 28920 28937 28948 29056
rect 28906 28928 28962 28937
rect 28906 28863 28962 28872
rect 29196 28257 29224 29514
rect 29276 29504 29328 29510
rect 29276 29446 29328 29452
rect 29288 29170 29316 29446
rect 29276 29164 29328 29170
rect 29276 29106 29328 29112
rect 29380 29102 29408 29786
rect 29460 29164 29512 29170
rect 29460 29106 29512 29112
rect 29368 29096 29420 29102
rect 29368 29038 29420 29044
rect 29472 28966 29500 29106
rect 29460 28960 29512 28966
rect 29460 28902 29512 28908
rect 29472 28558 29500 28902
rect 29460 28552 29512 28558
rect 29460 28494 29512 28500
rect 29564 28404 29592 31214
rect 29748 30938 29776 34886
rect 30208 34678 30236 34886
rect 30300 34678 30328 35022
rect 30196 34672 30248 34678
rect 30196 34614 30248 34620
rect 30288 34672 30340 34678
rect 30288 34614 30340 34620
rect 29828 34400 29880 34406
rect 29828 34342 29880 34348
rect 29840 33998 29868 34342
rect 30300 34202 30328 34614
rect 30392 34406 30420 35022
rect 30472 34944 30524 34950
rect 30472 34886 30524 34892
rect 30380 34400 30432 34406
rect 30380 34342 30432 34348
rect 29920 34196 29972 34202
rect 29920 34138 29972 34144
rect 30288 34196 30340 34202
rect 30288 34138 30340 34144
rect 29828 33992 29880 33998
rect 29828 33934 29880 33940
rect 29932 32910 29960 34138
rect 30288 33924 30340 33930
rect 30288 33866 30340 33872
rect 30196 33856 30248 33862
rect 30196 33798 30248 33804
rect 29920 32904 29972 32910
rect 29920 32846 29972 32852
rect 30208 32230 30236 33798
rect 30300 33658 30328 33866
rect 30288 33652 30340 33658
rect 30288 33594 30340 33600
rect 30392 32978 30420 34342
rect 30380 32972 30432 32978
rect 30380 32914 30432 32920
rect 30484 32502 30512 34886
rect 30748 33992 30800 33998
rect 30748 33934 30800 33940
rect 30656 32836 30708 32842
rect 30656 32778 30708 32784
rect 30472 32496 30524 32502
rect 30472 32438 30524 32444
rect 30380 32428 30432 32434
rect 30380 32370 30432 32376
rect 30196 32224 30248 32230
rect 30196 32166 30248 32172
rect 30208 31822 30236 32166
rect 30196 31816 30248 31822
rect 30196 31758 30248 31764
rect 29828 31340 29880 31346
rect 29828 31282 29880 31288
rect 29840 31210 29868 31282
rect 29828 31204 29880 31210
rect 29828 31146 29880 31152
rect 29736 30932 29788 30938
rect 29736 30874 29788 30880
rect 29748 30258 29776 30874
rect 29736 30252 29788 30258
rect 29736 30194 29788 30200
rect 29644 29096 29696 29102
rect 29644 29038 29696 29044
rect 29472 28376 29592 28404
rect 29182 28248 29238 28257
rect 29182 28183 29238 28192
rect 28724 28144 28776 28150
rect 28724 28086 28776 28092
rect 28816 28144 28868 28150
rect 28816 28086 28868 28092
rect 28920 28082 29132 28098
rect 28908 28076 29132 28082
rect 28960 28070 29132 28076
rect 28908 28018 28960 28024
rect 29104 28064 29132 28070
rect 29184 28076 29236 28082
rect 29104 28036 29184 28064
rect 29000 27872 29052 27878
rect 28998 27840 29000 27849
rect 29052 27840 29054 27849
rect 28998 27775 29054 27784
rect 28724 27600 28776 27606
rect 28724 27542 28776 27548
rect 28632 25832 28684 25838
rect 28632 25774 28684 25780
rect 28540 25696 28592 25702
rect 28540 25638 28592 25644
rect 28552 25294 28580 25638
rect 28644 25362 28672 25774
rect 28632 25356 28684 25362
rect 28632 25298 28684 25304
rect 28540 25288 28592 25294
rect 28540 25230 28592 25236
rect 28736 24188 28764 27542
rect 28816 26920 28868 26926
rect 28816 26862 28868 26868
rect 29000 26920 29052 26926
rect 29000 26862 29052 26868
rect 28828 26761 28856 26862
rect 28814 26752 28870 26761
rect 28814 26687 28870 26696
rect 28828 26314 28856 26687
rect 29012 26450 29040 26862
rect 29104 26790 29132 28036
rect 29368 28076 29420 28082
rect 29184 28018 29236 28024
rect 29288 28036 29368 28064
rect 29182 27976 29238 27985
rect 29182 27911 29238 27920
rect 29092 26784 29144 26790
rect 29092 26726 29144 26732
rect 29000 26444 29052 26450
rect 29000 26386 29052 26392
rect 28816 26308 28868 26314
rect 28816 26250 28868 26256
rect 29000 26308 29052 26314
rect 29000 26250 29052 26256
rect 28908 25968 28960 25974
rect 28908 25910 28960 25916
rect 28816 25832 28868 25838
rect 28816 25774 28868 25780
rect 28828 25430 28856 25774
rect 28816 25424 28868 25430
rect 28816 25366 28868 25372
rect 28920 24818 28948 25910
rect 28908 24812 28960 24818
rect 28908 24754 28960 24760
rect 28816 24200 28868 24206
rect 28736 24160 28816 24188
rect 28816 24142 28868 24148
rect 28540 24132 28592 24138
rect 28540 24074 28592 24080
rect 28552 23322 28580 24074
rect 28816 24064 28868 24070
rect 28816 24006 28868 24012
rect 28540 23316 28592 23322
rect 28540 23258 28592 23264
rect 28828 23118 28856 24006
rect 29012 23526 29040 26250
rect 29104 25974 29132 26726
rect 29196 26450 29224 27911
rect 29288 26772 29316 28036
rect 29368 28018 29420 28024
rect 29366 27976 29422 27985
rect 29366 27911 29422 27920
rect 29380 27470 29408 27911
rect 29368 27464 29420 27470
rect 29368 27406 29420 27412
rect 29472 26926 29500 28376
rect 29552 28212 29604 28218
rect 29552 28154 29604 28160
rect 29564 27690 29592 28154
rect 29656 28014 29684 29038
rect 29736 28960 29788 28966
rect 29736 28902 29788 28908
rect 29748 28082 29776 28902
rect 29736 28076 29788 28082
rect 29736 28018 29788 28024
rect 29644 28008 29696 28014
rect 29644 27950 29696 27956
rect 29644 27872 29696 27878
rect 29642 27840 29644 27849
rect 29696 27840 29698 27849
rect 29642 27775 29698 27784
rect 29642 27704 29698 27713
rect 29564 27662 29642 27690
rect 29642 27639 29698 27648
rect 29656 27470 29684 27639
rect 29644 27464 29696 27470
rect 29644 27406 29696 27412
rect 29736 27464 29788 27470
rect 29736 27406 29788 27412
rect 29748 27062 29776 27406
rect 29736 27056 29788 27062
rect 29736 26998 29788 27004
rect 29644 26988 29696 26994
rect 29644 26930 29696 26936
rect 29460 26920 29512 26926
rect 29460 26862 29512 26868
rect 29288 26744 29500 26772
rect 29656 26761 29684 26930
rect 29184 26444 29236 26450
rect 29184 26386 29236 26392
rect 29092 25968 29144 25974
rect 29092 25910 29144 25916
rect 29368 25968 29420 25974
rect 29368 25910 29420 25916
rect 29092 25220 29144 25226
rect 29092 25162 29144 25168
rect 29104 23866 29132 25162
rect 29276 24676 29328 24682
rect 29276 24618 29328 24624
rect 29092 23860 29144 23866
rect 29092 23802 29144 23808
rect 29288 23730 29316 24618
rect 29276 23724 29328 23730
rect 29276 23666 29328 23672
rect 29000 23520 29052 23526
rect 29000 23462 29052 23468
rect 29012 23304 29040 23462
rect 29012 23276 29132 23304
rect 29000 23180 29052 23186
rect 29000 23122 29052 23128
rect 28816 23112 28868 23118
rect 28816 23054 28868 23060
rect 28632 23044 28684 23050
rect 28632 22986 28684 22992
rect 28540 22636 28592 22642
rect 28540 22578 28592 22584
rect 28448 22228 28500 22234
rect 28448 22170 28500 22176
rect 28552 22166 28580 22578
rect 28540 22160 28592 22166
rect 28540 22102 28592 22108
rect 28264 22092 28316 22098
rect 28264 22034 28316 22040
rect 28552 21894 28580 22102
rect 28540 21888 28592 21894
rect 28540 21830 28592 21836
rect 28644 21690 28672 22986
rect 28724 22704 28776 22710
rect 28724 22646 28776 22652
rect 28736 22438 28764 22646
rect 29012 22574 29040 23122
rect 29104 22642 29132 23276
rect 29092 22636 29144 22642
rect 29092 22578 29144 22584
rect 29000 22568 29052 22574
rect 29000 22510 29052 22516
rect 29012 22438 29040 22510
rect 28724 22432 28776 22438
rect 28724 22374 28776 22380
rect 29000 22432 29052 22438
rect 29000 22374 29052 22380
rect 29012 22030 29040 22374
rect 29104 22094 29132 22578
rect 29104 22066 29224 22094
rect 29000 22024 29052 22030
rect 29000 21966 29052 21972
rect 28724 21888 28776 21894
rect 28724 21830 28776 21836
rect 28540 21684 28592 21690
rect 28540 21626 28592 21632
rect 28632 21684 28684 21690
rect 28632 21626 28684 21632
rect 28356 21344 28408 21350
rect 28356 21286 28408 21292
rect 28368 20942 28396 21286
rect 28448 21004 28500 21010
rect 28448 20946 28500 20952
rect 28356 20936 28408 20942
rect 28356 20878 28408 20884
rect 28368 20058 28396 20878
rect 28460 20874 28488 20946
rect 28552 20942 28580 21626
rect 28736 21554 28764 21830
rect 29000 21684 29052 21690
rect 29000 21626 29052 21632
rect 28724 21548 28776 21554
rect 28724 21490 28776 21496
rect 28908 21548 28960 21554
rect 28908 21490 28960 21496
rect 28920 20942 28948 21490
rect 28540 20936 28592 20942
rect 28540 20878 28592 20884
rect 28908 20936 28960 20942
rect 28908 20878 28960 20884
rect 28448 20868 28500 20874
rect 28448 20810 28500 20816
rect 28356 20052 28408 20058
rect 28356 19994 28408 20000
rect 28460 19854 28488 20810
rect 29012 20466 29040 21626
rect 29092 21616 29144 21622
rect 29092 21558 29144 21564
rect 28632 20460 28684 20466
rect 28632 20402 28684 20408
rect 29000 20460 29052 20466
rect 29000 20402 29052 20408
rect 28448 19848 28500 19854
rect 28448 19790 28500 19796
rect 28172 19712 28224 19718
rect 28172 19654 28224 19660
rect 28448 19712 28500 19718
rect 28448 19654 28500 19660
rect 28460 19378 28488 19654
rect 28448 19372 28500 19378
rect 28448 19314 28500 19320
rect 28644 18154 28672 20402
rect 28724 20392 28776 20398
rect 28724 20334 28776 20340
rect 28736 20058 28764 20334
rect 28724 20052 28776 20058
rect 28724 19994 28776 20000
rect 29012 19854 29040 20402
rect 29000 19848 29052 19854
rect 29000 19790 29052 19796
rect 28908 19780 28960 19786
rect 28908 19722 28960 19728
rect 28920 19689 28948 19722
rect 28906 19680 28962 19689
rect 28906 19615 28962 19624
rect 29012 19378 29040 19790
rect 29000 19372 29052 19378
rect 29000 19314 29052 19320
rect 28722 19272 28778 19281
rect 28722 19207 28724 19216
rect 28776 19207 28778 19216
rect 28724 19178 28776 19184
rect 29104 19174 29132 21558
rect 29196 21554 29224 22066
rect 29184 21548 29236 21554
rect 29184 21490 29236 21496
rect 29288 20942 29316 23666
rect 29380 23361 29408 25910
rect 29472 25294 29500 26744
rect 29642 26752 29698 26761
rect 29642 26687 29698 26696
rect 29460 25288 29512 25294
rect 29460 25230 29512 25236
rect 29366 23352 29422 23361
rect 29366 23287 29422 23296
rect 29368 23180 29420 23186
rect 29368 23122 29420 23128
rect 29380 22642 29408 23122
rect 29368 22636 29420 22642
rect 29368 22578 29420 22584
rect 29368 21548 29420 21554
rect 29368 21490 29420 21496
rect 29276 20936 29328 20942
rect 29276 20878 29328 20884
rect 29184 20800 29236 20806
rect 29184 20742 29236 20748
rect 29196 20534 29224 20742
rect 29184 20528 29236 20534
rect 29184 20470 29236 20476
rect 29196 20330 29224 20470
rect 29184 20324 29236 20330
rect 29184 20266 29236 20272
rect 29288 20074 29316 20878
rect 29380 20806 29408 21490
rect 29368 20800 29420 20806
rect 29368 20742 29420 20748
rect 29196 20046 29316 20074
rect 29092 19168 29144 19174
rect 29092 19110 29144 19116
rect 28724 18624 28776 18630
rect 28724 18566 28776 18572
rect 28736 18290 28764 18566
rect 28724 18284 28776 18290
rect 28724 18226 28776 18232
rect 28632 18148 28684 18154
rect 28632 18090 28684 18096
rect 29196 18086 29224 20046
rect 29276 19984 29328 19990
rect 29276 19926 29328 19932
rect 29288 18970 29316 19926
rect 29380 19854 29408 20742
rect 29368 19848 29420 19854
rect 29368 19790 29420 19796
rect 29368 19168 29420 19174
rect 29368 19110 29420 19116
rect 29276 18964 29328 18970
rect 29276 18906 29328 18912
rect 29380 18902 29408 19110
rect 29368 18896 29420 18902
rect 29368 18838 29420 18844
rect 29472 18766 29500 25230
rect 29656 24206 29684 26687
rect 29736 25900 29788 25906
rect 29736 25842 29788 25848
rect 29644 24200 29696 24206
rect 29644 24142 29696 24148
rect 29644 24064 29696 24070
rect 29644 24006 29696 24012
rect 29656 23798 29684 24006
rect 29644 23792 29696 23798
rect 29644 23734 29696 23740
rect 29644 23656 29696 23662
rect 29644 23598 29696 23604
rect 29552 22024 29604 22030
rect 29552 21966 29604 21972
rect 29564 21418 29592 21966
rect 29656 21690 29684 23598
rect 29644 21684 29696 21690
rect 29644 21626 29696 21632
rect 29552 21412 29604 21418
rect 29552 21354 29604 21360
rect 29644 21344 29696 21350
rect 29644 21286 29696 21292
rect 29656 21010 29684 21286
rect 29644 21004 29696 21010
rect 29644 20946 29696 20952
rect 29748 19854 29776 25842
rect 29840 23798 29868 31146
rect 30104 31136 30156 31142
rect 30104 31078 30156 31084
rect 30116 30870 30144 31078
rect 30392 30938 30420 32370
rect 30484 31414 30512 32438
rect 30564 32360 30616 32366
rect 30564 32302 30616 32308
rect 30576 31890 30604 32302
rect 30564 31884 30616 31890
rect 30564 31826 30616 31832
rect 30576 31793 30604 31826
rect 30562 31784 30618 31793
rect 30562 31719 30618 31728
rect 30564 31476 30616 31482
rect 30564 31418 30616 31424
rect 30472 31408 30524 31414
rect 30472 31350 30524 31356
rect 30472 31272 30524 31278
rect 30472 31214 30524 31220
rect 30484 31142 30512 31214
rect 30472 31136 30524 31142
rect 30472 31078 30524 31084
rect 30380 30932 30432 30938
rect 30380 30874 30432 30880
rect 30104 30864 30156 30870
rect 30104 30806 30156 30812
rect 30288 30592 30340 30598
rect 30288 30534 30340 30540
rect 30300 30190 30328 30534
rect 30380 30388 30432 30394
rect 30380 30330 30432 30336
rect 29920 30184 29972 30190
rect 29920 30126 29972 30132
rect 30288 30184 30340 30190
rect 30288 30126 30340 30132
rect 29932 29510 29960 30126
rect 30012 29572 30064 29578
rect 30012 29514 30064 29520
rect 29920 29504 29972 29510
rect 29920 29446 29972 29452
rect 29932 25702 29960 29446
rect 30024 29306 30052 29514
rect 30104 29504 30156 29510
rect 30104 29446 30156 29452
rect 30012 29300 30064 29306
rect 30012 29242 30064 29248
rect 30024 27441 30052 29242
rect 30116 29102 30144 29446
rect 30104 29096 30156 29102
rect 30104 29038 30156 29044
rect 30104 28960 30156 28966
rect 30104 28902 30156 28908
rect 30116 28014 30144 28902
rect 30196 28416 30248 28422
rect 30196 28358 30248 28364
rect 30104 28008 30156 28014
rect 30104 27950 30156 27956
rect 30010 27432 30066 27441
rect 30010 27367 30066 27376
rect 30104 27056 30156 27062
rect 30104 26998 30156 27004
rect 30012 26988 30064 26994
rect 30012 26930 30064 26936
rect 30024 26382 30052 26930
rect 30116 26625 30144 26998
rect 30102 26616 30158 26625
rect 30102 26551 30158 26560
rect 30012 26376 30064 26382
rect 30010 26344 30012 26353
rect 30064 26344 30066 26353
rect 30010 26279 30066 26288
rect 30024 26253 30052 26279
rect 30012 26036 30064 26042
rect 30012 25978 30064 25984
rect 29920 25696 29972 25702
rect 29920 25638 29972 25644
rect 30024 25362 30052 25978
rect 30208 25922 30236 28358
rect 30300 28014 30328 30126
rect 30392 29170 30420 30330
rect 30484 30190 30512 31078
rect 30472 30184 30524 30190
rect 30472 30126 30524 30132
rect 30576 30002 30604 31418
rect 30484 29974 30604 30002
rect 30380 29164 30432 29170
rect 30380 29106 30432 29112
rect 30392 28762 30420 29106
rect 30380 28756 30432 28762
rect 30380 28698 30432 28704
rect 30380 28552 30432 28558
rect 30380 28494 30432 28500
rect 30288 28008 30340 28014
rect 30288 27950 30340 27956
rect 30392 27470 30420 28494
rect 30484 27470 30512 29974
rect 30668 29866 30696 32778
rect 30760 32774 30788 33934
rect 30840 33856 30892 33862
rect 30840 33798 30892 33804
rect 30748 32768 30800 32774
rect 30748 32710 30800 32716
rect 30760 31929 30788 32710
rect 30746 31920 30802 31929
rect 30746 31855 30802 31864
rect 30746 31512 30802 31521
rect 30746 31447 30802 31456
rect 30576 29838 30696 29866
rect 30576 29034 30604 29838
rect 30656 29708 30708 29714
rect 30656 29650 30708 29656
rect 30668 29170 30696 29650
rect 30656 29164 30708 29170
rect 30656 29106 30708 29112
rect 30564 29028 30616 29034
rect 30564 28970 30616 28976
rect 30564 28688 30616 28694
rect 30564 28630 30616 28636
rect 30380 27464 30432 27470
rect 30380 27406 30432 27412
rect 30472 27464 30524 27470
rect 30472 27406 30524 27412
rect 30380 27328 30432 27334
rect 30380 27270 30432 27276
rect 30472 27328 30524 27334
rect 30472 27270 30524 27276
rect 30392 26432 30420 27270
rect 30116 25906 30236 25922
rect 30300 26404 30420 26432
rect 30300 25906 30328 26404
rect 30484 26382 30512 27270
rect 30576 26994 30604 28630
rect 30760 27538 30788 31447
rect 30852 29730 30880 33798
rect 30944 32978 30972 35090
rect 31024 34604 31076 34610
rect 31024 34546 31076 34552
rect 31036 34406 31064 34546
rect 31024 34400 31076 34406
rect 31024 34342 31076 34348
rect 31220 33980 31248 36110
rect 31300 36100 31352 36106
rect 31300 36042 31352 36048
rect 31312 35698 31340 36042
rect 31300 35692 31352 35698
rect 31300 35634 31352 35640
rect 31300 35488 31352 35494
rect 31300 35430 31352 35436
rect 31312 34048 31340 35430
rect 31588 35086 31616 36314
rect 32128 36236 32180 36242
rect 32128 36178 32180 36184
rect 31668 36168 31720 36174
rect 31668 36110 31720 36116
rect 31680 35290 31708 36110
rect 31852 36032 31904 36038
rect 31852 35974 31904 35980
rect 31864 35630 31892 35974
rect 32140 35698 32168 36178
rect 32220 36168 32272 36174
rect 32220 36110 32272 36116
rect 32404 36168 32456 36174
rect 32404 36110 32456 36116
rect 32128 35692 32180 35698
rect 32128 35634 32180 35640
rect 31852 35624 31904 35630
rect 31852 35566 31904 35572
rect 32140 35290 32168 35634
rect 32232 35630 32260 36110
rect 32220 35624 32272 35630
rect 32220 35566 32272 35572
rect 32416 35578 32444 36110
rect 32508 35834 32536 36586
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 32956 36032 33008 36038
rect 32956 35974 33008 35980
rect 32496 35828 32548 35834
rect 32496 35770 32548 35776
rect 32968 35698 32996 35974
rect 32956 35692 33008 35698
rect 32956 35634 33008 35640
rect 31668 35284 31720 35290
rect 31668 35226 31720 35232
rect 32128 35284 32180 35290
rect 32128 35226 32180 35232
rect 31680 35086 31708 35226
rect 31576 35080 31628 35086
rect 31576 35022 31628 35028
rect 31668 35080 31720 35086
rect 31668 35022 31720 35028
rect 31392 34944 31444 34950
rect 31392 34886 31444 34892
rect 31404 34746 31432 34886
rect 31392 34740 31444 34746
rect 31392 34682 31444 34688
rect 31588 34678 31616 35022
rect 31576 34672 31628 34678
rect 31576 34614 31628 34620
rect 32232 34610 32260 35566
rect 32416 35550 32536 35578
rect 32508 35494 32536 35550
rect 32496 35488 32548 35494
rect 32496 35430 32548 35436
rect 33048 35488 33100 35494
rect 33048 35430 33100 35436
rect 32220 34604 32272 34610
rect 32220 34546 32272 34552
rect 31392 34400 31444 34406
rect 31392 34342 31444 34348
rect 31760 34400 31812 34406
rect 31760 34342 31812 34348
rect 31404 34202 31432 34342
rect 31392 34196 31444 34202
rect 31392 34138 31444 34144
rect 31668 34128 31720 34134
rect 31668 34070 31720 34076
rect 31312 34020 31432 34048
rect 31220 33952 31340 33980
rect 31208 33856 31260 33862
rect 31208 33798 31260 33804
rect 31220 33590 31248 33798
rect 31208 33584 31260 33590
rect 31208 33526 31260 33532
rect 31312 33522 31340 33952
rect 31404 33522 31432 34020
rect 31680 33862 31708 34070
rect 31668 33856 31720 33862
rect 31668 33798 31720 33804
rect 31668 33584 31720 33590
rect 31668 33526 31720 33532
rect 31300 33516 31352 33522
rect 31300 33458 31352 33464
rect 31392 33516 31444 33522
rect 31392 33458 31444 33464
rect 31300 33312 31352 33318
rect 31300 33254 31352 33260
rect 31208 33040 31260 33046
rect 31208 32982 31260 32988
rect 30932 32972 30984 32978
rect 30932 32914 30984 32920
rect 30944 32366 30972 32914
rect 30932 32360 30984 32366
rect 30932 32302 30984 32308
rect 31024 32292 31076 32298
rect 31024 32234 31076 32240
rect 30930 32056 30986 32065
rect 30930 31991 30986 32000
rect 30944 31890 30972 31991
rect 30932 31884 30984 31890
rect 30932 31826 30984 31832
rect 30944 31346 30972 31826
rect 30932 31340 30984 31346
rect 30932 31282 30984 31288
rect 31036 30938 31064 32234
rect 31116 32224 31168 32230
rect 31116 32166 31168 32172
rect 31024 30932 31076 30938
rect 31024 30874 31076 30880
rect 31128 30734 31156 32166
rect 31220 31210 31248 32982
rect 31312 32434 31340 33254
rect 31404 32502 31432 33458
rect 31484 32836 31536 32842
rect 31484 32778 31536 32784
rect 31392 32496 31444 32502
rect 31392 32438 31444 32444
rect 31496 32434 31524 32778
rect 31680 32570 31708 33526
rect 31772 33046 31800 34342
rect 31944 34128 31996 34134
rect 31944 34070 31996 34076
rect 31956 33998 31984 34070
rect 31944 33992 31996 33998
rect 31944 33934 31996 33940
rect 31956 33522 31984 33934
rect 32232 33930 32260 34546
rect 32404 34536 32456 34542
rect 32404 34478 32456 34484
rect 32312 34400 32364 34406
rect 32312 34342 32364 34348
rect 32220 33924 32272 33930
rect 32220 33866 32272 33872
rect 31944 33516 31996 33522
rect 31944 33458 31996 33464
rect 32324 33454 32352 34342
rect 32416 34066 32444 34478
rect 32404 34060 32456 34066
rect 32404 34002 32456 34008
rect 32312 33448 32364 33454
rect 32312 33390 32364 33396
rect 31852 33380 31904 33386
rect 31852 33322 31904 33328
rect 31760 33040 31812 33046
rect 31760 32982 31812 32988
rect 31864 32910 31892 33322
rect 32508 33114 32536 35430
rect 33060 35222 33088 35430
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 33048 35216 33100 35222
rect 33048 35158 33100 35164
rect 34612 34672 34664 34678
rect 34612 34614 34664 34620
rect 33048 34060 33100 34066
rect 33048 34002 33100 34008
rect 32772 33992 32824 33998
rect 32772 33934 32824 33940
rect 32680 33924 32732 33930
rect 32680 33866 32732 33872
rect 32588 33312 32640 33318
rect 32588 33254 32640 33260
rect 32496 33108 32548 33114
rect 32496 33050 32548 33056
rect 31852 32904 31904 32910
rect 31852 32846 31904 32852
rect 32496 32904 32548 32910
rect 32496 32846 32548 32852
rect 31760 32836 31812 32842
rect 31760 32778 31812 32784
rect 31576 32564 31628 32570
rect 31576 32506 31628 32512
rect 31668 32564 31720 32570
rect 31668 32506 31720 32512
rect 31588 32450 31616 32506
rect 31300 32428 31352 32434
rect 31300 32370 31352 32376
rect 31484 32428 31536 32434
rect 31588 32422 31708 32450
rect 31484 32370 31536 32376
rect 31312 31804 31340 32370
rect 31496 32298 31524 32370
rect 31576 32360 31628 32366
rect 31576 32302 31628 32308
rect 31484 32292 31536 32298
rect 31484 32234 31536 32240
rect 31496 32065 31524 32234
rect 31482 32056 31538 32065
rect 31482 31991 31538 32000
rect 31588 31958 31616 32302
rect 31576 31952 31628 31958
rect 31576 31894 31628 31900
rect 31392 31816 31444 31822
rect 31312 31776 31392 31804
rect 31392 31758 31444 31764
rect 31484 31748 31536 31754
rect 31484 31690 31536 31696
rect 31300 31408 31352 31414
rect 31300 31350 31352 31356
rect 31208 31204 31260 31210
rect 31208 31146 31260 31152
rect 31116 30728 31168 30734
rect 31116 30670 31168 30676
rect 30932 30660 30984 30666
rect 30932 30602 30984 30608
rect 30944 30054 30972 30602
rect 31312 30394 31340 31350
rect 31496 31226 31524 31690
rect 31576 31680 31628 31686
rect 31576 31622 31628 31628
rect 31404 31198 31524 31226
rect 31404 30666 31432 31198
rect 31484 31136 31536 31142
rect 31484 31078 31536 31084
rect 31496 30938 31524 31078
rect 31588 30938 31616 31622
rect 31680 31142 31708 32422
rect 31772 32366 31800 32778
rect 31760 32360 31812 32366
rect 31760 32302 31812 32308
rect 31760 32224 31812 32230
rect 31760 32166 31812 32172
rect 31668 31136 31720 31142
rect 31668 31078 31720 31084
rect 31772 30954 31800 32166
rect 31864 31754 31892 32846
rect 31944 32836 31996 32842
rect 31944 32778 31996 32784
rect 31852 31748 31904 31754
rect 31852 31690 31904 31696
rect 31864 31346 31892 31690
rect 31852 31340 31904 31346
rect 31852 31282 31904 31288
rect 31484 30932 31536 30938
rect 31484 30874 31536 30880
rect 31576 30932 31628 30938
rect 31576 30874 31628 30880
rect 31680 30926 31800 30954
rect 31588 30802 31616 30874
rect 31576 30796 31628 30802
rect 31576 30738 31628 30744
rect 31392 30660 31444 30666
rect 31392 30602 31444 30608
rect 31300 30388 31352 30394
rect 31300 30330 31352 30336
rect 30932 30048 30984 30054
rect 30932 29990 30984 29996
rect 30852 29702 31616 29730
rect 31208 29640 31260 29646
rect 31208 29582 31260 29588
rect 31220 29170 31248 29582
rect 31208 29164 31260 29170
rect 31260 29124 31340 29152
rect 31208 29106 31260 29112
rect 31208 29028 31260 29034
rect 31208 28970 31260 28976
rect 31024 28756 31076 28762
rect 31024 28698 31076 28704
rect 30930 28656 30986 28665
rect 30930 28591 30986 28600
rect 30944 28218 30972 28591
rect 31036 28558 31064 28698
rect 31024 28552 31076 28558
rect 31024 28494 31076 28500
rect 31114 28384 31170 28393
rect 31114 28319 31170 28328
rect 30932 28212 30984 28218
rect 30932 28154 30984 28160
rect 31128 28150 31156 28319
rect 31116 28144 31168 28150
rect 31116 28086 31168 28092
rect 30840 28076 30892 28082
rect 30840 28018 30892 28024
rect 30932 28076 30984 28082
rect 30932 28018 30984 28024
rect 30852 27849 30880 28018
rect 30838 27840 30894 27849
rect 30838 27775 30894 27784
rect 30748 27532 30800 27538
rect 30748 27474 30800 27480
rect 30656 27464 30708 27470
rect 30656 27406 30708 27412
rect 30840 27464 30892 27470
rect 30840 27406 30892 27412
rect 30668 27010 30696 27406
rect 30564 26988 30616 26994
rect 30668 26982 30788 27010
rect 30852 26994 30880 27406
rect 30564 26930 30616 26936
rect 30656 26920 30708 26926
rect 30656 26862 30708 26868
rect 30564 26784 30616 26790
rect 30564 26726 30616 26732
rect 30472 26376 30524 26382
rect 30472 26318 30524 26324
rect 30380 26308 30432 26314
rect 30380 26250 30432 26256
rect 30104 25900 30236 25906
rect 30156 25894 30236 25900
rect 30288 25900 30340 25906
rect 30104 25842 30156 25848
rect 30288 25842 30340 25848
rect 30300 25702 30328 25842
rect 30288 25696 30340 25702
rect 30288 25638 30340 25644
rect 30392 25514 30420 26250
rect 30392 25486 30512 25514
rect 30380 25424 30432 25430
rect 30380 25366 30432 25372
rect 30012 25356 30064 25362
rect 30012 25298 30064 25304
rect 30392 24750 30420 25366
rect 30380 24744 30432 24750
rect 30380 24686 30432 24692
rect 29828 23792 29880 23798
rect 29828 23734 29880 23740
rect 29840 22166 29868 23734
rect 30392 23186 30420 24686
rect 30380 23180 30432 23186
rect 30380 23122 30432 23128
rect 30484 22642 30512 25486
rect 30472 22636 30524 22642
rect 30472 22578 30524 22584
rect 29920 22432 29972 22438
rect 29920 22374 29972 22380
rect 29828 22160 29880 22166
rect 29828 22102 29880 22108
rect 29840 22030 29868 22102
rect 29828 22024 29880 22030
rect 29828 21966 29880 21972
rect 29932 21622 29960 22374
rect 30576 22234 30604 26726
rect 30668 26518 30696 26862
rect 30656 26512 30708 26518
rect 30656 26454 30708 26460
rect 30668 26382 30696 26454
rect 30656 26376 30708 26382
rect 30656 26318 30708 26324
rect 30760 25786 30788 26982
rect 30840 26988 30892 26994
rect 30840 26930 30892 26936
rect 30852 25906 30880 26930
rect 30944 26330 30972 28018
rect 31128 27606 31156 28086
rect 31116 27600 31168 27606
rect 31116 27542 31168 27548
rect 31024 27532 31076 27538
rect 31024 27474 31076 27480
rect 31036 26450 31064 27474
rect 31220 27452 31248 28970
rect 31128 27424 31248 27452
rect 31024 26444 31076 26450
rect 31024 26386 31076 26392
rect 30944 26302 31064 26330
rect 30930 26208 30986 26217
rect 30930 26143 30986 26152
rect 30944 25974 30972 26143
rect 30932 25968 30984 25974
rect 30932 25910 30984 25916
rect 30840 25900 30892 25906
rect 30840 25842 30892 25848
rect 30656 25764 30708 25770
rect 30760 25758 30880 25786
rect 30656 25706 30708 25712
rect 30668 25294 30696 25706
rect 30748 25696 30800 25702
rect 30748 25638 30800 25644
rect 30656 25288 30708 25294
rect 30656 25230 30708 25236
rect 30760 25158 30788 25638
rect 30656 25152 30708 25158
rect 30656 25094 30708 25100
rect 30748 25152 30800 25158
rect 30748 25094 30800 25100
rect 30668 24818 30696 25094
rect 30746 24984 30802 24993
rect 30746 24919 30802 24928
rect 30656 24812 30708 24818
rect 30656 24754 30708 24760
rect 30656 24200 30708 24206
rect 30656 24142 30708 24148
rect 30668 23662 30696 24142
rect 30760 23730 30788 24919
rect 30852 24410 30880 25758
rect 30944 25265 30972 25910
rect 31036 25906 31064 26302
rect 31024 25900 31076 25906
rect 31024 25842 31076 25848
rect 31024 25492 31076 25498
rect 31024 25434 31076 25440
rect 30930 25256 30986 25265
rect 30930 25191 30986 25200
rect 30932 25152 30984 25158
rect 30932 25094 30984 25100
rect 30840 24404 30892 24410
rect 30840 24346 30892 24352
rect 30748 23724 30800 23730
rect 30748 23666 30800 23672
rect 30656 23656 30708 23662
rect 30656 23598 30708 23604
rect 30668 22574 30696 23598
rect 30852 23050 30880 24346
rect 30840 23044 30892 23050
rect 30840 22986 30892 22992
rect 30656 22568 30708 22574
rect 30656 22510 30708 22516
rect 30564 22228 30616 22234
rect 30564 22170 30616 22176
rect 30748 22092 30800 22098
rect 30748 22034 30800 22040
rect 30656 21956 30708 21962
rect 30656 21898 30708 21904
rect 30012 21888 30064 21894
rect 30012 21830 30064 21836
rect 30104 21888 30156 21894
rect 30104 21830 30156 21836
rect 30024 21690 30052 21830
rect 30012 21684 30064 21690
rect 30012 21626 30064 21632
rect 29920 21616 29972 21622
rect 29920 21558 29972 21564
rect 29920 20596 29972 20602
rect 29920 20538 29972 20544
rect 29736 19848 29788 19854
rect 29736 19790 29788 19796
rect 29552 19712 29604 19718
rect 29552 19654 29604 19660
rect 29564 19378 29592 19654
rect 29932 19514 29960 20538
rect 30116 20534 30144 21830
rect 30668 21604 30696 21898
rect 30760 21729 30788 22034
rect 30840 21888 30892 21894
rect 30840 21830 30892 21836
rect 30746 21720 30802 21729
rect 30746 21655 30802 21664
rect 30852 21604 30880 21830
rect 30562 21584 30618 21593
rect 30668 21576 30880 21604
rect 30562 21519 30618 21528
rect 30576 21486 30604 21519
rect 30564 21480 30616 21486
rect 30564 21422 30616 21428
rect 30748 21412 30800 21418
rect 30748 21354 30800 21360
rect 30564 21344 30616 21350
rect 30564 21286 30616 21292
rect 30104 20528 30156 20534
rect 30104 20470 30156 20476
rect 30576 19854 30604 21286
rect 30760 20874 30788 21354
rect 30748 20868 30800 20874
rect 30748 20810 30800 20816
rect 30564 19848 30616 19854
rect 30564 19790 30616 19796
rect 30472 19712 30524 19718
rect 30472 19654 30524 19660
rect 29920 19508 29972 19514
rect 29920 19450 29972 19456
rect 29644 19440 29696 19446
rect 29642 19408 29644 19417
rect 29696 19408 29698 19417
rect 29552 19372 29604 19378
rect 29642 19343 29698 19352
rect 29552 19314 29604 19320
rect 29932 18766 29960 19450
rect 30378 19408 30434 19417
rect 30378 19343 30434 19352
rect 30196 19304 30248 19310
rect 30196 19246 30248 19252
rect 30208 18766 30236 19246
rect 29460 18760 29512 18766
rect 29460 18702 29512 18708
rect 29736 18760 29788 18766
rect 29736 18702 29788 18708
rect 29920 18760 29972 18766
rect 29920 18702 29972 18708
rect 30196 18760 30248 18766
rect 30196 18702 30248 18708
rect 29748 18426 29776 18702
rect 30104 18692 30156 18698
rect 30104 18634 30156 18640
rect 29736 18420 29788 18426
rect 29736 18362 29788 18368
rect 27988 18080 28040 18086
rect 27988 18022 28040 18028
rect 29184 18080 29236 18086
rect 29184 18022 29236 18028
rect 30116 17882 30144 18634
rect 30208 18358 30236 18702
rect 30196 18352 30248 18358
rect 30196 18294 30248 18300
rect 30392 17882 30420 19343
rect 30484 18970 30512 19654
rect 30576 19446 30604 19790
rect 30564 19440 30616 19446
rect 30564 19382 30616 19388
rect 30472 18964 30524 18970
rect 30472 18906 30524 18912
rect 30852 18766 30880 21576
rect 30944 21554 30972 25094
rect 31036 24886 31064 25434
rect 31024 24880 31076 24886
rect 31024 24822 31076 24828
rect 31036 24206 31064 24822
rect 31024 24200 31076 24206
rect 31024 24142 31076 24148
rect 31036 22982 31064 24142
rect 31024 22976 31076 22982
rect 31024 22918 31076 22924
rect 31024 22772 31076 22778
rect 31024 22714 31076 22720
rect 30932 21548 30984 21554
rect 30932 21490 30984 21496
rect 31036 21010 31064 22714
rect 31024 21004 31076 21010
rect 31024 20946 31076 20952
rect 30932 20936 30984 20942
rect 30932 20878 30984 20884
rect 30944 20602 30972 20878
rect 30932 20596 30984 20602
rect 30932 20538 30984 20544
rect 31128 19854 31156 27424
rect 31312 26024 31340 29124
rect 31484 28620 31536 28626
rect 31484 28562 31536 28568
rect 31496 28218 31524 28562
rect 31484 28212 31536 28218
rect 31484 28154 31536 28160
rect 31392 28008 31444 28014
rect 31392 27950 31444 27956
rect 31404 27033 31432 27950
rect 31482 27568 31538 27577
rect 31482 27503 31538 27512
rect 31496 27470 31524 27503
rect 31484 27464 31536 27470
rect 31484 27406 31536 27412
rect 31484 27328 31536 27334
rect 31482 27296 31484 27305
rect 31536 27296 31538 27305
rect 31482 27231 31538 27240
rect 31390 27024 31446 27033
rect 31390 26959 31446 26968
rect 31588 26926 31616 29702
rect 31392 26920 31444 26926
rect 31392 26862 31444 26868
rect 31576 26920 31628 26926
rect 31576 26862 31628 26868
rect 31220 25996 31340 26024
rect 31220 25498 31248 25996
rect 31300 25900 31352 25906
rect 31300 25842 31352 25848
rect 31208 25492 31260 25498
rect 31208 25434 31260 25440
rect 31208 25288 31260 25294
rect 31208 25230 31260 25236
rect 31220 24750 31248 25230
rect 31312 25226 31340 25842
rect 31404 25838 31432 26862
rect 31484 26784 31536 26790
rect 31484 26726 31536 26732
rect 31392 25832 31444 25838
rect 31392 25774 31444 25780
rect 31392 25696 31444 25702
rect 31392 25638 31444 25644
rect 31300 25220 31352 25226
rect 31300 25162 31352 25168
rect 31404 25106 31432 25638
rect 31312 25078 31432 25106
rect 31312 24886 31340 25078
rect 31300 24880 31352 24886
rect 31300 24822 31352 24828
rect 31208 24744 31260 24750
rect 31208 24686 31260 24692
rect 31208 24064 31260 24070
rect 31208 24006 31260 24012
rect 31220 22030 31248 24006
rect 31208 22024 31260 22030
rect 31208 21966 31260 21972
rect 31220 21418 31248 21966
rect 31312 21554 31340 24822
rect 31496 23322 31524 26726
rect 31576 26512 31628 26518
rect 31576 26454 31628 26460
rect 31588 24954 31616 26454
rect 31680 25922 31708 30926
rect 31852 30864 31904 30870
rect 31852 30806 31904 30812
rect 31864 29714 31892 30806
rect 31956 30258 31984 32778
rect 32508 32570 32536 32846
rect 32496 32564 32548 32570
rect 32496 32506 32548 32512
rect 32220 32428 32272 32434
rect 32220 32370 32272 32376
rect 32312 32428 32364 32434
rect 32312 32370 32364 32376
rect 32232 31822 32260 32370
rect 32324 31822 32352 32370
rect 32600 31958 32628 33254
rect 32692 32910 32720 33866
rect 32784 33590 32812 33934
rect 32772 33584 32824 33590
rect 32772 33526 32824 33532
rect 32680 32904 32732 32910
rect 32680 32846 32732 32852
rect 32692 32502 32720 32846
rect 32784 32842 32812 33526
rect 32864 33516 32916 33522
rect 32864 33458 32916 33464
rect 32876 32910 32904 33458
rect 33060 32978 33088 34002
rect 33876 33992 33928 33998
rect 33876 33934 33928 33940
rect 33888 33454 33916 33934
rect 33876 33448 33928 33454
rect 33876 33390 33928 33396
rect 33416 33040 33468 33046
rect 33416 32982 33468 32988
rect 33048 32972 33100 32978
rect 33048 32914 33100 32920
rect 32864 32904 32916 32910
rect 32864 32846 32916 32852
rect 32956 32904 33008 32910
rect 32956 32846 33008 32852
rect 32772 32836 32824 32842
rect 32772 32778 32824 32784
rect 32680 32496 32732 32502
rect 32680 32438 32732 32444
rect 32968 32026 32996 32846
rect 33324 32224 33376 32230
rect 33324 32166 33376 32172
rect 32956 32020 33008 32026
rect 32956 31962 33008 31968
rect 32588 31952 32640 31958
rect 32588 31894 32640 31900
rect 32600 31822 32628 31894
rect 32968 31822 32996 31962
rect 33048 31884 33100 31890
rect 33048 31826 33100 31832
rect 33232 31884 33284 31890
rect 33232 31826 33284 31832
rect 32220 31816 32272 31822
rect 32220 31758 32272 31764
rect 32312 31816 32364 31822
rect 32312 31758 32364 31764
rect 32588 31816 32640 31822
rect 32588 31758 32640 31764
rect 32956 31816 33008 31822
rect 32956 31758 33008 31764
rect 33060 31770 33088 31826
rect 33060 31742 33180 31770
rect 32036 31680 32088 31686
rect 32036 31622 32088 31628
rect 32048 31278 32076 31622
rect 33152 31482 33180 31742
rect 33140 31476 33192 31482
rect 33140 31418 33192 31424
rect 32128 31340 32180 31346
rect 32128 31282 32180 31288
rect 32036 31272 32088 31278
rect 32036 31214 32088 31220
rect 32140 30598 32168 31282
rect 32588 31272 32640 31278
rect 32588 31214 32640 31220
rect 32864 31272 32916 31278
rect 32864 31214 32916 31220
rect 32600 30734 32628 31214
rect 32680 31136 32732 31142
rect 32680 31078 32732 31084
rect 32692 30938 32720 31078
rect 32680 30932 32732 30938
rect 32680 30874 32732 30880
rect 32588 30728 32640 30734
rect 32588 30670 32640 30676
rect 32772 30660 32824 30666
rect 32772 30602 32824 30608
rect 32128 30592 32180 30598
rect 32128 30534 32180 30540
rect 32220 30320 32272 30326
rect 32140 30268 32220 30274
rect 32272 30268 32536 30274
rect 32140 30258 32536 30268
rect 31944 30252 31996 30258
rect 31944 30194 31996 30200
rect 32140 30252 32548 30258
rect 32140 30246 32496 30252
rect 31852 29708 31904 29714
rect 31852 29650 31904 29656
rect 31864 28966 31892 29650
rect 31956 29306 31984 30194
rect 31944 29300 31996 29306
rect 31944 29242 31996 29248
rect 32036 29232 32088 29238
rect 32036 29174 32088 29180
rect 31852 28960 31904 28966
rect 31852 28902 31904 28908
rect 31852 28620 31904 28626
rect 31852 28562 31904 28568
rect 31864 28490 31892 28562
rect 32048 28558 32076 29174
rect 32036 28552 32088 28558
rect 32034 28520 32036 28529
rect 32088 28520 32090 28529
rect 31852 28484 31904 28490
rect 32034 28455 32090 28464
rect 31852 28426 31904 28432
rect 32140 28370 32168 30246
rect 32496 30194 32548 30200
rect 32312 30048 32364 30054
rect 32312 29990 32364 29996
rect 32220 29708 32272 29714
rect 32220 29650 32272 29656
rect 32232 29510 32260 29650
rect 32220 29504 32272 29510
rect 32220 29446 32272 29452
rect 32232 28694 32260 29446
rect 32324 29306 32352 29990
rect 32496 29640 32548 29646
rect 32496 29582 32548 29588
rect 32312 29300 32364 29306
rect 32312 29242 32364 29248
rect 32220 28688 32272 28694
rect 32220 28630 32272 28636
rect 32232 28558 32260 28630
rect 32220 28552 32272 28558
rect 32220 28494 32272 28500
rect 32324 28490 32352 29242
rect 32508 28994 32536 29582
rect 32680 29300 32732 29306
rect 32680 29242 32732 29248
rect 32692 29034 32720 29242
rect 32416 28966 32536 28994
rect 32680 29028 32732 29034
rect 32680 28970 32732 28976
rect 32312 28484 32364 28490
rect 32312 28426 32364 28432
rect 32048 28342 32168 28370
rect 32220 28416 32272 28422
rect 32220 28358 32272 28364
rect 31852 28144 31904 28150
rect 31850 28112 31852 28121
rect 31904 28112 31906 28121
rect 31772 28070 31850 28098
rect 31772 27402 31800 28070
rect 31850 28047 31906 28056
rect 31944 28076 31996 28082
rect 31944 28018 31996 28024
rect 31956 27878 31984 28018
rect 32048 27946 32076 28342
rect 32126 28248 32182 28257
rect 32126 28183 32182 28192
rect 32036 27940 32088 27946
rect 32036 27882 32088 27888
rect 31944 27872 31996 27878
rect 31996 27820 32076 27826
rect 31944 27814 32076 27820
rect 31956 27798 32076 27814
rect 31942 27704 31998 27713
rect 31942 27639 31944 27648
rect 31996 27639 31998 27648
rect 31944 27610 31996 27616
rect 31852 27600 31904 27606
rect 31850 27568 31852 27577
rect 31904 27568 31906 27577
rect 32048 27538 32076 27798
rect 31850 27503 31906 27512
rect 31944 27532 31996 27538
rect 31944 27474 31996 27480
rect 32036 27532 32088 27538
rect 32036 27474 32088 27480
rect 31852 27464 31904 27470
rect 31852 27406 31904 27412
rect 31760 27396 31812 27402
rect 31760 27338 31812 27344
rect 31864 27305 31892 27406
rect 31850 27296 31906 27305
rect 31850 27231 31906 27240
rect 31760 26920 31812 26926
rect 31760 26862 31812 26868
rect 31772 26586 31800 26862
rect 31852 26852 31904 26858
rect 31852 26794 31904 26800
rect 31760 26580 31812 26586
rect 31760 26522 31812 26528
rect 31864 26314 31892 26794
rect 31956 26450 31984 27474
rect 32034 27024 32090 27033
rect 32034 26959 32090 26968
rect 31944 26444 31996 26450
rect 31944 26386 31996 26392
rect 31852 26308 31904 26314
rect 31852 26250 31904 26256
rect 31956 25974 31984 26386
rect 32048 26042 32076 26959
rect 32036 26036 32088 26042
rect 32036 25978 32088 25984
rect 31944 25968 31996 25974
rect 31680 25894 31800 25922
rect 31944 25910 31996 25916
rect 31668 25764 31720 25770
rect 31668 25706 31720 25712
rect 31680 25378 31708 25706
rect 31772 25514 31800 25894
rect 31772 25486 31892 25514
rect 31680 25350 31800 25378
rect 31576 24948 31628 24954
rect 31576 24890 31628 24896
rect 31576 24608 31628 24614
rect 31772 24596 31800 25350
rect 31864 24614 31892 25486
rect 31944 24948 31996 24954
rect 31944 24890 31996 24896
rect 31576 24550 31628 24556
rect 31680 24568 31800 24596
rect 31852 24608 31904 24614
rect 31484 23316 31536 23322
rect 31404 23276 31484 23304
rect 31404 22642 31432 23276
rect 31484 23258 31536 23264
rect 31484 23112 31536 23118
rect 31484 23054 31536 23060
rect 31392 22636 31444 22642
rect 31392 22578 31444 22584
rect 31496 22574 31524 23054
rect 31484 22568 31536 22574
rect 31484 22510 31536 22516
rect 31588 22098 31616 24550
rect 31576 22092 31628 22098
rect 31576 22034 31628 22040
rect 31576 21616 31628 21622
rect 31576 21558 31628 21564
rect 31300 21548 31352 21554
rect 31300 21490 31352 21496
rect 31208 21412 31260 21418
rect 31208 21354 31260 21360
rect 31588 21010 31616 21558
rect 31576 21004 31628 21010
rect 31576 20946 31628 20952
rect 31680 20806 31708 24568
rect 31852 24550 31904 24556
rect 31956 23186 31984 24890
rect 32048 24818 32076 25978
rect 32036 24812 32088 24818
rect 32036 24754 32088 24760
rect 32036 24676 32088 24682
rect 32036 24618 32088 24624
rect 32048 23798 32076 24618
rect 32036 23792 32088 23798
rect 32036 23734 32088 23740
rect 32140 23254 32168 28183
rect 32232 27713 32260 28358
rect 32416 28150 32444 28966
rect 32680 28416 32732 28422
rect 32680 28358 32732 28364
rect 32692 28257 32720 28358
rect 32678 28248 32734 28257
rect 32678 28183 32734 28192
rect 32404 28144 32456 28150
rect 32324 28104 32404 28132
rect 32218 27704 32274 27713
rect 32218 27639 32274 27648
rect 32324 27632 32352 28104
rect 32404 28086 32456 28092
rect 32784 28082 32812 30602
rect 32876 29714 32904 31214
rect 32956 30320 33008 30326
rect 32956 30262 33008 30268
rect 32864 29708 32916 29714
rect 32864 29650 32916 29656
rect 32772 28076 32824 28082
rect 32772 28018 32824 28024
rect 32404 27940 32456 27946
rect 32404 27882 32456 27888
rect 32680 27940 32732 27946
rect 32680 27882 32732 27888
rect 32416 27632 32444 27882
rect 32586 27840 32642 27849
rect 32586 27775 32642 27784
rect 32496 27668 32548 27674
rect 32312 27626 32364 27632
rect 32312 27568 32364 27574
rect 32404 27626 32456 27632
rect 32496 27610 32548 27616
rect 32404 27568 32456 27574
rect 32508 27452 32536 27610
rect 32416 27441 32536 27452
rect 32402 27432 32536 27441
rect 32458 27424 32536 27432
rect 32402 27367 32458 27376
rect 32416 26994 32444 27367
rect 32496 27056 32548 27062
rect 32496 26998 32548 27004
rect 32220 26988 32272 26994
rect 32404 26988 32456 26994
rect 32272 26948 32404 26976
rect 32220 26930 32272 26936
rect 32404 26930 32456 26936
rect 32508 26897 32536 26998
rect 32494 26888 32550 26897
rect 32494 26823 32550 26832
rect 32508 26382 32536 26823
rect 32600 26450 32628 27775
rect 32588 26444 32640 26450
rect 32588 26386 32640 26392
rect 32496 26376 32548 26382
rect 32496 26318 32548 26324
rect 32508 26042 32536 26318
rect 32496 26036 32548 26042
rect 32496 25978 32548 25984
rect 32312 25900 32364 25906
rect 32312 25842 32364 25848
rect 32324 25294 32352 25842
rect 32496 25696 32548 25702
rect 32496 25638 32548 25644
rect 32312 25288 32364 25294
rect 32312 25230 32364 25236
rect 32220 25152 32272 25158
rect 32220 25094 32272 25100
rect 32232 24206 32260 25094
rect 32404 24608 32456 24614
rect 32404 24550 32456 24556
rect 32220 24200 32272 24206
rect 32220 24142 32272 24148
rect 32312 24200 32364 24206
rect 32312 24142 32364 24148
rect 32128 23248 32180 23254
rect 32128 23190 32180 23196
rect 31944 23180 31996 23186
rect 31944 23122 31996 23128
rect 31956 22710 31984 23122
rect 31944 22704 31996 22710
rect 31944 22646 31996 22652
rect 32128 22500 32180 22506
rect 32128 22442 32180 22448
rect 32140 21554 32168 22442
rect 32232 22030 32260 24142
rect 32324 23866 32352 24142
rect 32416 24070 32444 24550
rect 32508 24274 32536 25638
rect 32692 24342 32720 27882
rect 32876 26625 32904 29650
rect 32968 29510 32996 30262
rect 33048 30252 33100 30258
rect 33048 30194 33100 30200
rect 32956 29504 33008 29510
rect 32956 29446 33008 29452
rect 32968 29170 32996 29446
rect 33060 29306 33088 30194
rect 33244 29866 33272 31826
rect 33336 30870 33364 32166
rect 33428 31822 33456 32982
rect 33784 32768 33836 32774
rect 33784 32710 33836 32716
rect 33796 32570 33824 32710
rect 33784 32564 33836 32570
rect 33784 32506 33836 32512
rect 33888 32502 33916 33390
rect 33968 32904 34020 32910
rect 33968 32846 34020 32852
rect 33508 32496 33560 32502
rect 33508 32438 33560 32444
rect 33876 32496 33928 32502
rect 33876 32438 33928 32444
rect 33520 32026 33548 32438
rect 33508 32020 33560 32026
rect 33508 31962 33560 31968
rect 33416 31816 33468 31822
rect 33416 31758 33468 31764
rect 33980 30938 34008 32846
rect 34152 31952 34204 31958
rect 34152 31894 34204 31900
rect 34164 31822 34192 31894
rect 34152 31816 34204 31822
rect 34152 31758 34204 31764
rect 34060 31748 34112 31754
rect 34060 31690 34112 31696
rect 33968 30932 34020 30938
rect 33968 30874 34020 30880
rect 33324 30864 33376 30870
rect 33324 30806 33376 30812
rect 33600 30728 33652 30734
rect 33600 30670 33652 30676
rect 33244 29838 33548 29866
rect 33232 29708 33284 29714
rect 33232 29650 33284 29656
rect 33244 29306 33272 29650
rect 33048 29300 33100 29306
rect 33048 29242 33100 29248
rect 33232 29300 33284 29306
rect 33232 29242 33284 29248
rect 32956 29164 33008 29170
rect 32956 29106 33008 29112
rect 33232 29096 33284 29102
rect 33232 29038 33284 29044
rect 33048 28960 33100 28966
rect 33048 28902 33100 28908
rect 32954 28384 33010 28393
rect 32954 28319 33010 28328
rect 32862 26616 32918 26625
rect 32862 26551 32918 26560
rect 32772 26376 32824 26382
rect 32772 26318 32824 26324
rect 32784 25974 32812 26318
rect 32772 25968 32824 25974
rect 32772 25910 32824 25916
rect 32876 25294 32904 26551
rect 32968 25906 32996 28319
rect 33060 27878 33088 28902
rect 33244 28121 33272 29038
rect 33416 28620 33468 28626
rect 33416 28562 33468 28568
rect 33428 28393 33456 28562
rect 33414 28384 33470 28393
rect 33414 28319 33470 28328
rect 33230 28112 33286 28121
rect 33230 28047 33286 28056
rect 33048 27872 33100 27878
rect 33048 27814 33100 27820
rect 33232 27464 33284 27470
rect 33232 27406 33284 27412
rect 33048 27124 33100 27130
rect 33048 27066 33100 27072
rect 33140 27124 33192 27130
rect 33140 27066 33192 27072
rect 33060 26858 33088 27066
rect 33048 26852 33100 26858
rect 33048 26794 33100 26800
rect 33048 26240 33100 26246
rect 33152 26194 33180 27066
rect 33244 26790 33272 27406
rect 33416 27328 33468 27334
rect 33322 27296 33378 27305
rect 33416 27270 33468 27276
rect 33322 27231 33378 27240
rect 33336 27062 33364 27231
rect 33324 27056 33376 27062
rect 33324 26998 33376 27004
rect 33232 26784 33284 26790
rect 33232 26726 33284 26732
rect 33244 26314 33272 26726
rect 33428 26586 33456 27270
rect 33520 26926 33548 29838
rect 33612 29782 33640 30670
rect 34072 30666 34100 31690
rect 34520 31680 34572 31686
rect 34520 31622 34572 31628
rect 34532 31346 34560 31622
rect 34520 31340 34572 31346
rect 34520 31282 34572 31288
rect 34624 31278 34652 34614
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 34796 33380 34848 33386
rect 34796 33322 34848 33328
rect 34808 32978 34836 33322
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 34796 32972 34848 32978
rect 34796 32914 34848 32920
rect 34704 32292 34756 32298
rect 34704 32234 34756 32240
rect 34716 31958 34744 32234
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 35624 32020 35676 32026
rect 35624 31962 35676 31968
rect 34704 31952 34756 31958
rect 34704 31894 34756 31900
rect 34716 31822 34744 31894
rect 35532 31884 35584 31890
rect 35532 31826 35584 31832
rect 34704 31816 34756 31822
rect 34704 31758 34756 31764
rect 35544 31346 35572 31826
rect 35636 31754 35664 31962
rect 35636 31726 35756 31754
rect 35532 31340 35584 31346
rect 35532 31282 35584 31288
rect 34612 31272 34664 31278
rect 34612 31214 34664 31220
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 35072 30728 35124 30734
rect 35072 30670 35124 30676
rect 35624 30728 35676 30734
rect 35624 30670 35676 30676
rect 34060 30660 34112 30666
rect 34060 30602 34112 30608
rect 33968 30048 34020 30054
rect 33968 29990 34020 29996
rect 33600 29776 33652 29782
rect 33600 29718 33652 29724
rect 33980 29646 34008 29990
rect 33968 29640 34020 29646
rect 33968 29582 34020 29588
rect 33784 29572 33836 29578
rect 33784 29514 33836 29520
rect 33796 28762 33824 29514
rect 33876 29164 33928 29170
rect 33876 29106 33928 29112
rect 33784 28756 33836 28762
rect 33784 28698 33836 28704
rect 33888 28490 33916 29106
rect 33968 29096 34020 29102
rect 33968 29038 34020 29044
rect 33980 28665 34008 29038
rect 33966 28656 34022 28665
rect 33966 28591 34022 28600
rect 33980 28558 34008 28591
rect 33968 28552 34020 28558
rect 33968 28494 34020 28500
rect 33876 28484 33928 28490
rect 33876 28426 33928 28432
rect 33600 28144 33652 28150
rect 33600 28086 33652 28092
rect 33612 27418 33640 28086
rect 33692 28076 33744 28082
rect 33692 28018 33744 28024
rect 33704 27985 33732 28018
rect 33968 28008 34020 28014
rect 33690 27976 33746 27985
rect 33968 27950 34020 27956
rect 33690 27911 33746 27920
rect 33876 27872 33928 27878
rect 33876 27814 33928 27820
rect 33612 27390 33824 27418
rect 33508 26920 33560 26926
rect 33508 26862 33560 26868
rect 33416 26580 33468 26586
rect 33416 26522 33468 26528
rect 33612 26489 33640 27390
rect 33796 27334 33824 27390
rect 33692 27328 33744 27334
rect 33692 27270 33744 27276
rect 33784 27328 33836 27334
rect 33784 27270 33836 27276
rect 33704 27062 33732 27270
rect 33888 27130 33916 27814
rect 33876 27124 33928 27130
rect 33876 27066 33928 27072
rect 33692 27056 33744 27062
rect 33692 26998 33744 27004
rect 33598 26480 33654 26489
rect 33598 26415 33654 26424
rect 33508 26376 33560 26382
rect 33508 26318 33560 26324
rect 33232 26308 33284 26314
rect 33232 26250 33284 26256
rect 33100 26188 33180 26194
rect 33048 26182 33180 26188
rect 33060 26166 33180 26182
rect 33152 25906 33180 26166
rect 32956 25900 33008 25906
rect 32956 25842 33008 25848
rect 33140 25900 33192 25906
rect 33140 25842 33192 25848
rect 32864 25288 32916 25294
rect 32864 25230 32916 25236
rect 33152 24886 33180 25842
rect 33140 24880 33192 24886
rect 33140 24822 33192 24828
rect 32772 24812 32824 24818
rect 32772 24754 32824 24760
rect 32784 24682 32812 24754
rect 32772 24676 32824 24682
rect 32772 24618 32824 24624
rect 32680 24336 32732 24342
rect 32680 24278 32732 24284
rect 32496 24268 32548 24274
rect 32496 24210 32548 24216
rect 32404 24064 32456 24070
rect 32404 24006 32456 24012
rect 32312 23860 32364 23866
rect 32312 23802 32364 23808
rect 32692 23730 32720 24278
rect 33152 24274 33180 24822
rect 33140 24268 33192 24274
rect 33140 24210 33192 24216
rect 32956 24064 33008 24070
rect 32956 24006 33008 24012
rect 32680 23724 32732 23730
rect 32680 23666 32732 23672
rect 32968 23050 32996 24006
rect 33048 23724 33100 23730
rect 33048 23666 33100 23672
rect 33060 23322 33088 23666
rect 33152 23662 33180 24210
rect 33244 24206 33272 26250
rect 33520 26246 33548 26318
rect 33508 26240 33560 26246
rect 33508 26182 33560 26188
rect 33520 25974 33548 26182
rect 33508 25968 33560 25974
rect 33508 25910 33560 25916
rect 33704 25158 33732 26998
rect 33782 26752 33838 26761
rect 33782 26687 33838 26696
rect 33796 26042 33824 26687
rect 33876 26444 33928 26450
rect 33980 26432 34008 27950
rect 34072 26450 34100 30602
rect 35084 30394 35112 30670
rect 35072 30388 35124 30394
rect 35072 30330 35124 30336
rect 35636 30326 35664 30670
rect 35624 30320 35676 30326
rect 35624 30262 35676 30268
rect 34152 30252 34204 30258
rect 34152 30194 34204 30200
rect 34164 29782 34192 30194
rect 34796 30116 34848 30122
rect 34796 30058 34848 30064
rect 34704 29844 34756 29850
rect 34704 29786 34756 29792
rect 34152 29776 34204 29782
rect 34152 29718 34204 29724
rect 34716 29646 34744 29786
rect 34808 29714 34836 30058
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 34796 29708 34848 29714
rect 34796 29650 34848 29656
rect 34520 29640 34572 29646
rect 34520 29582 34572 29588
rect 34704 29640 34756 29646
rect 34704 29582 34756 29588
rect 34336 29300 34388 29306
rect 34336 29242 34388 29248
rect 34150 29200 34206 29209
rect 34150 29135 34206 29144
rect 34164 29034 34192 29135
rect 34152 29028 34204 29034
rect 34152 28970 34204 28976
rect 34348 28694 34376 29242
rect 34532 29102 34560 29582
rect 34808 29238 34836 29650
rect 35636 29646 35664 30262
rect 34980 29640 35032 29646
rect 34980 29582 35032 29588
rect 35624 29640 35676 29646
rect 35624 29582 35676 29588
rect 34888 29504 34940 29510
rect 34888 29446 34940 29452
rect 34796 29232 34848 29238
rect 34796 29174 34848 29180
rect 34900 29170 34928 29446
rect 34992 29306 35020 29582
rect 34980 29300 35032 29306
rect 34980 29242 35032 29248
rect 34704 29164 34756 29170
rect 34704 29106 34756 29112
rect 34888 29164 34940 29170
rect 34888 29106 34940 29112
rect 34520 29096 34572 29102
rect 34520 29038 34572 29044
rect 34428 28960 34480 28966
rect 34428 28902 34480 28908
rect 34336 28688 34388 28694
rect 34336 28630 34388 28636
rect 34440 28218 34468 28902
rect 34532 28558 34560 29038
rect 34612 29028 34664 29034
rect 34612 28970 34664 28976
rect 34520 28552 34572 28558
rect 34520 28494 34572 28500
rect 34428 28212 34480 28218
rect 34428 28154 34480 28160
rect 34520 28076 34572 28082
rect 34520 28018 34572 28024
rect 34532 27674 34560 28018
rect 34520 27668 34572 27674
rect 34520 27610 34572 27616
rect 34624 27554 34652 28970
rect 34716 28694 34744 29106
rect 35532 29096 35584 29102
rect 35532 29038 35584 29044
rect 34796 28960 34848 28966
rect 34796 28902 34848 28908
rect 34704 28688 34756 28694
rect 34704 28630 34756 28636
rect 34808 28626 34836 28902
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 35544 28762 35572 29038
rect 35532 28756 35584 28762
rect 35532 28698 35584 28704
rect 34796 28620 34848 28626
rect 34796 28562 34848 28568
rect 35440 28076 35492 28082
rect 35440 28018 35492 28024
rect 34794 27976 34850 27985
rect 34794 27911 34850 27920
rect 34428 27532 34480 27538
rect 34624 27526 34744 27554
rect 34428 27474 34480 27480
rect 34440 26926 34468 27474
rect 34612 27464 34664 27470
rect 34612 27406 34664 27412
rect 34624 26994 34652 27406
rect 34612 26988 34664 26994
rect 34612 26930 34664 26936
rect 34428 26920 34480 26926
rect 34428 26862 34480 26868
rect 34520 26852 34572 26858
rect 34520 26794 34572 26800
rect 34532 26518 34560 26794
rect 34336 26512 34388 26518
rect 34336 26454 34388 26460
rect 34520 26512 34572 26518
rect 34520 26454 34572 26460
rect 33928 26404 34008 26432
rect 34060 26444 34112 26450
rect 33876 26386 33928 26392
rect 34060 26386 34112 26392
rect 34072 26353 34100 26386
rect 34058 26344 34114 26353
rect 34058 26279 34114 26288
rect 33784 26036 33836 26042
rect 33784 25978 33836 25984
rect 34348 25906 34376 26454
rect 34624 26314 34652 26930
rect 34612 26308 34664 26314
rect 34612 26250 34664 26256
rect 34336 25900 34388 25906
rect 34336 25842 34388 25848
rect 33876 25696 33928 25702
rect 33876 25638 33928 25644
rect 33692 25152 33744 25158
rect 33692 25094 33744 25100
rect 33704 24732 33732 25094
rect 33888 24818 33916 25638
rect 34060 25356 34112 25362
rect 34060 25298 34112 25304
rect 34072 24954 34100 25298
rect 34060 24948 34112 24954
rect 34060 24890 34112 24896
rect 34348 24818 34376 25842
rect 34520 25696 34572 25702
rect 34520 25638 34572 25644
rect 34532 25362 34560 25638
rect 34716 25378 34744 27526
rect 34808 26382 34836 27911
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 35072 27328 35124 27334
rect 35072 27270 35124 27276
rect 35084 26994 35112 27270
rect 35072 26988 35124 26994
rect 35072 26930 35124 26936
rect 35348 26784 35400 26790
rect 35348 26726 35400 26732
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 35360 26625 35388 26726
rect 35346 26616 35402 26625
rect 35346 26551 35402 26560
rect 34980 26512 35032 26518
rect 34980 26454 35032 26460
rect 34992 26382 35020 26454
rect 34796 26376 34848 26382
rect 34796 26318 34848 26324
rect 34980 26376 35032 26382
rect 34980 26318 35032 26324
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 34796 25492 34848 25498
rect 34796 25434 34848 25440
rect 34520 25356 34572 25362
rect 34520 25298 34572 25304
rect 34624 25350 34744 25378
rect 33876 24812 33928 24818
rect 33876 24754 33928 24760
rect 34336 24812 34388 24818
rect 34336 24754 34388 24760
rect 33784 24744 33836 24750
rect 33704 24704 33784 24732
rect 33784 24686 33836 24692
rect 33232 24200 33284 24206
rect 33232 24142 33284 24148
rect 33692 23860 33744 23866
rect 33692 23802 33744 23808
rect 33600 23724 33652 23730
rect 33600 23666 33652 23672
rect 33140 23656 33192 23662
rect 33140 23598 33192 23604
rect 33140 23520 33192 23526
rect 33140 23462 33192 23468
rect 33048 23316 33100 23322
rect 33048 23258 33100 23264
rect 33152 23118 33180 23462
rect 33140 23112 33192 23118
rect 33140 23054 33192 23060
rect 32956 23044 33008 23050
rect 32956 22986 33008 22992
rect 32864 22636 32916 22642
rect 32968 22624 32996 22986
rect 33152 22778 33180 23054
rect 33232 22976 33284 22982
rect 33232 22918 33284 22924
rect 33416 22976 33468 22982
rect 33416 22918 33468 22924
rect 33140 22772 33192 22778
rect 33140 22714 33192 22720
rect 32916 22596 32996 22624
rect 32864 22578 32916 22584
rect 33244 22574 33272 22918
rect 33232 22568 33284 22574
rect 33232 22510 33284 22516
rect 33232 22432 33284 22438
rect 33232 22374 33284 22380
rect 32496 22092 32548 22098
rect 32496 22034 32548 22040
rect 32220 22024 32272 22030
rect 32220 21966 32272 21972
rect 32508 21894 32536 22034
rect 32496 21888 32548 21894
rect 32496 21830 32548 21836
rect 32508 21690 32536 21830
rect 32496 21684 32548 21690
rect 32496 21626 32548 21632
rect 32128 21548 32180 21554
rect 32128 21490 32180 21496
rect 32140 20942 32168 21490
rect 32404 21344 32456 21350
rect 32404 21286 32456 21292
rect 32416 20942 32444 21286
rect 33048 21072 33100 21078
rect 33048 21014 33100 21020
rect 32128 20936 32180 20942
rect 32128 20878 32180 20884
rect 32404 20936 32456 20942
rect 32404 20878 32456 20884
rect 32496 20868 32548 20874
rect 32496 20810 32548 20816
rect 31668 20800 31720 20806
rect 31668 20742 31720 20748
rect 32036 20800 32088 20806
rect 32036 20742 32088 20748
rect 32048 20466 32076 20742
rect 32508 20466 32536 20810
rect 32036 20460 32088 20466
rect 32036 20402 32088 20408
rect 32128 20460 32180 20466
rect 32128 20402 32180 20408
rect 32496 20460 32548 20466
rect 32496 20402 32548 20408
rect 31668 20392 31720 20398
rect 31668 20334 31720 20340
rect 31680 19854 31708 20334
rect 31760 20256 31812 20262
rect 31760 20198 31812 20204
rect 31116 19848 31168 19854
rect 31116 19790 31168 19796
rect 31668 19848 31720 19854
rect 31668 19790 31720 19796
rect 31024 19712 31076 19718
rect 31024 19654 31076 19660
rect 31036 18766 31064 19654
rect 31128 19446 31156 19790
rect 31116 19440 31168 19446
rect 31116 19382 31168 19388
rect 31772 19310 31800 20198
rect 32048 19922 32076 20402
rect 32140 20058 32168 20402
rect 32588 20256 32640 20262
rect 32588 20198 32640 20204
rect 32772 20256 32824 20262
rect 32772 20198 32824 20204
rect 32128 20052 32180 20058
rect 32128 19994 32180 20000
rect 32036 19916 32088 19922
rect 32036 19858 32088 19864
rect 32140 19378 32168 19994
rect 32404 19712 32456 19718
rect 32404 19654 32456 19660
rect 32128 19372 32180 19378
rect 32128 19314 32180 19320
rect 31760 19304 31812 19310
rect 31760 19246 31812 19252
rect 31116 19168 31168 19174
rect 31116 19110 31168 19116
rect 31300 19168 31352 19174
rect 31300 19110 31352 19116
rect 30840 18760 30892 18766
rect 30840 18702 30892 18708
rect 31024 18760 31076 18766
rect 31024 18702 31076 18708
rect 30104 17876 30156 17882
rect 30104 17818 30156 17824
rect 30380 17876 30432 17882
rect 30380 17818 30432 17824
rect 30852 17678 30880 18702
rect 30840 17672 30892 17678
rect 30840 17614 30892 17620
rect 31036 17542 31064 18702
rect 31128 18630 31156 19110
rect 31116 18624 31168 18630
rect 31116 18566 31168 18572
rect 31128 18222 31156 18566
rect 31208 18420 31260 18426
rect 31208 18362 31260 18368
rect 31116 18216 31168 18222
rect 31116 18158 31168 18164
rect 31220 17814 31248 18362
rect 31312 18290 31340 19110
rect 31772 18970 31800 19246
rect 31760 18964 31812 18970
rect 31760 18906 31812 18912
rect 31668 18760 31720 18766
rect 31668 18702 31720 18708
rect 31392 18352 31444 18358
rect 31392 18294 31444 18300
rect 31300 18284 31352 18290
rect 31300 18226 31352 18232
rect 31404 17882 31432 18294
rect 31680 18290 31708 18702
rect 31668 18284 31720 18290
rect 31668 18226 31720 18232
rect 31484 18216 31536 18222
rect 31484 18158 31536 18164
rect 31392 17876 31444 17882
rect 31392 17818 31444 17824
rect 31208 17808 31260 17814
rect 31208 17750 31260 17756
rect 31496 17678 31524 18158
rect 31772 18086 31800 18906
rect 31852 18760 31904 18766
rect 31852 18702 31904 18708
rect 31760 18080 31812 18086
rect 31760 18022 31812 18028
rect 31484 17672 31536 17678
rect 31484 17614 31536 17620
rect 31864 17610 31892 18702
rect 32140 18290 32168 19314
rect 32416 19242 32444 19654
rect 32600 19446 32628 20198
rect 32784 20058 32812 20198
rect 32772 20052 32824 20058
rect 32772 19994 32824 20000
rect 33060 19718 33088 21014
rect 33244 20942 33272 22374
rect 33428 22166 33456 22918
rect 33612 22710 33640 23666
rect 33704 23118 33732 23802
rect 34624 23662 34652 25350
rect 34808 24970 34836 25434
rect 35256 25288 35308 25294
rect 35256 25230 35308 25236
rect 34716 24942 34836 24970
rect 34716 24206 34744 24942
rect 35268 24886 35296 25230
rect 35256 24880 35308 24886
rect 35256 24822 35308 24828
rect 34796 24676 34848 24682
rect 34796 24618 34848 24624
rect 34808 24206 34836 24618
rect 35452 24614 35480 28018
rect 35624 27464 35676 27470
rect 35624 27406 35676 27412
rect 35636 27062 35664 27406
rect 35728 27169 35756 31726
rect 35714 27160 35770 27169
rect 35714 27095 35770 27104
rect 35624 27056 35676 27062
rect 35544 27004 35624 27010
rect 35544 26998 35676 27004
rect 35544 26982 35664 26998
rect 35728 26994 35756 27095
rect 35716 26988 35768 26994
rect 35544 26382 35572 26982
rect 35716 26930 35768 26936
rect 35624 26920 35676 26926
rect 35624 26862 35676 26868
rect 35636 26450 35664 26862
rect 35624 26444 35676 26450
rect 35624 26386 35676 26392
rect 35532 26376 35584 26382
rect 35532 26318 35584 26324
rect 35716 25968 35768 25974
rect 35716 25910 35768 25916
rect 35728 25226 35756 25910
rect 35716 25220 35768 25226
rect 35716 25162 35768 25168
rect 35440 24608 35492 24614
rect 35440 24550 35492 24556
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 34704 24200 34756 24206
rect 34704 24142 34756 24148
rect 34796 24200 34848 24206
rect 34796 24142 34848 24148
rect 35348 24200 35400 24206
rect 35348 24142 35400 24148
rect 34796 24064 34848 24070
rect 34796 24006 34848 24012
rect 34612 23656 34664 23662
rect 34612 23598 34664 23604
rect 34518 23216 34574 23225
rect 34518 23151 34574 23160
rect 33692 23112 33744 23118
rect 33692 23054 33744 23060
rect 33600 22704 33652 22710
rect 33600 22646 33652 22652
rect 33612 22506 33640 22646
rect 33600 22500 33652 22506
rect 33600 22442 33652 22448
rect 33704 22166 33732 23054
rect 33784 22976 33836 22982
rect 33784 22918 33836 22924
rect 33796 22166 33824 22918
rect 33968 22432 34020 22438
rect 33968 22374 34020 22380
rect 34428 22432 34480 22438
rect 34428 22374 34480 22380
rect 33416 22160 33468 22166
rect 33416 22102 33468 22108
rect 33692 22160 33744 22166
rect 33692 22102 33744 22108
rect 33784 22160 33836 22166
rect 33784 22102 33836 22108
rect 33980 21622 34008 22374
rect 34060 22024 34112 22030
rect 34060 21966 34112 21972
rect 34072 21690 34100 21966
rect 34060 21684 34112 21690
rect 34060 21626 34112 21632
rect 33968 21616 34020 21622
rect 33968 21558 34020 21564
rect 34440 21554 34468 22374
rect 34428 21548 34480 21554
rect 34428 21490 34480 21496
rect 33324 21140 33376 21146
rect 33324 21082 33376 21088
rect 33232 20936 33284 20942
rect 33232 20878 33284 20884
rect 33140 20800 33192 20806
rect 33140 20742 33192 20748
rect 33048 19712 33100 19718
rect 33048 19654 33100 19660
rect 32588 19440 32640 19446
rect 32588 19382 32640 19388
rect 32864 19440 32916 19446
rect 32864 19382 32916 19388
rect 32680 19372 32732 19378
rect 32680 19314 32732 19320
rect 32404 19236 32456 19242
rect 32404 19178 32456 19184
rect 32692 18766 32720 19314
rect 32876 18766 32904 19382
rect 33152 19242 33180 20742
rect 33244 20534 33272 20878
rect 33232 20528 33284 20534
rect 33232 20470 33284 20476
rect 33336 20398 33364 21082
rect 33876 20528 33928 20534
rect 33876 20470 33928 20476
rect 33324 20392 33376 20398
rect 33324 20334 33376 20340
rect 33888 19514 33916 20470
rect 34244 20256 34296 20262
rect 34244 20198 34296 20204
rect 34256 19922 34284 20198
rect 34244 19916 34296 19922
rect 34244 19858 34296 19864
rect 34336 19780 34388 19786
rect 34336 19722 34388 19728
rect 33876 19508 33928 19514
rect 33876 19450 33928 19456
rect 34060 19372 34112 19378
rect 34060 19314 34112 19320
rect 34152 19372 34204 19378
rect 34152 19314 34204 19320
rect 33140 19236 33192 19242
rect 33140 19178 33192 19184
rect 33152 18766 33180 19178
rect 33968 19168 34020 19174
rect 33968 19110 34020 19116
rect 33980 18766 34008 19110
rect 34072 18902 34100 19314
rect 34060 18896 34112 18902
rect 34060 18838 34112 18844
rect 32680 18760 32732 18766
rect 32680 18702 32732 18708
rect 32864 18760 32916 18766
rect 32864 18702 32916 18708
rect 33140 18760 33192 18766
rect 33140 18702 33192 18708
rect 33968 18760 34020 18766
rect 33968 18702 34020 18708
rect 32404 18624 32456 18630
rect 32404 18566 32456 18572
rect 32416 18358 32444 18566
rect 32692 18426 32720 18702
rect 33232 18692 33284 18698
rect 33232 18634 33284 18640
rect 32956 18624 33008 18630
rect 32956 18566 33008 18572
rect 32680 18420 32732 18426
rect 32680 18362 32732 18368
rect 32404 18352 32456 18358
rect 32404 18294 32456 18300
rect 32128 18284 32180 18290
rect 32128 18226 32180 18232
rect 32416 17678 32444 18294
rect 32968 18290 32996 18566
rect 33244 18426 33272 18634
rect 33980 18426 34008 18702
rect 33232 18420 33284 18426
rect 33232 18362 33284 18368
rect 33968 18420 34020 18426
rect 33968 18362 34020 18368
rect 32956 18284 33008 18290
rect 32956 18226 33008 18232
rect 32968 17746 32996 18226
rect 34072 18222 34100 18838
rect 34164 18290 34192 19314
rect 34152 18284 34204 18290
rect 34152 18226 34204 18232
rect 34348 18222 34376 19722
rect 34532 18834 34560 23151
rect 34808 23050 34836 24006
rect 35360 23866 35388 24142
rect 35624 24064 35676 24070
rect 35624 24006 35676 24012
rect 35348 23860 35400 23866
rect 35348 23802 35400 23808
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 35360 23118 35388 23802
rect 35636 23662 35664 24006
rect 35716 23860 35768 23866
rect 35716 23802 35768 23808
rect 35624 23656 35676 23662
rect 35624 23598 35676 23604
rect 35636 23322 35664 23598
rect 35624 23316 35676 23322
rect 35624 23258 35676 23264
rect 35348 23112 35400 23118
rect 35348 23054 35400 23060
rect 34796 23044 34848 23050
rect 34796 22986 34848 22992
rect 35440 22976 35492 22982
rect 35440 22918 35492 22924
rect 35636 22930 35664 23258
rect 35728 23050 35756 23802
rect 35716 23044 35768 23050
rect 35716 22986 35768 22992
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 34612 22228 34664 22234
rect 34612 22170 34664 22176
rect 34624 21622 34652 22170
rect 35452 22030 35480 22918
rect 35636 22902 35756 22930
rect 35624 22704 35676 22710
rect 35624 22646 35676 22652
rect 35532 22432 35584 22438
rect 35532 22374 35584 22380
rect 35440 22024 35492 22030
rect 35440 21966 35492 21972
rect 34704 21888 34756 21894
rect 34704 21830 34756 21836
rect 34716 21622 34744 21830
rect 34612 21616 34664 21622
rect 34612 21558 34664 21564
rect 34704 21616 34756 21622
rect 34704 21558 34756 21564
rect 35544 21554 35572 22374
rect 35636 22234 35664 22646
rect 35624 22228 35676 22234
rect 35624 22170 35676 22176
rect 35728 22094 35756 22902
rect 35636 22066 35756 22094
rect 35636 22030 35664 22066
rect 35624 22024 35676 22030
rect 35624 21966 35676 21972
rect 35532 21548 35584 21554
rect 35532 21490 35584 21496
rect 34796 21344 34848 21350
rect 34796 21286 34848 21292
rect 34612 21004 34664 21010
rect 34612 20946 34664 20952
rect 34624 19378 34652 20946
rect 34704 20936 34756 20942
rect 34704 20878 34756 20884
rect 34716 20466 34744 20878
rect 34808 20534 34836 21286
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 34888 21072 34940 21078
rect 34888 21014 34940 21020
rect 34900 20874 34928 21014
rect 35544 20942 35572 21490
rect 35716 21480 35768 21486
rect 35716 21422 35768 21428
rect 35624 21072 35676 21078
rect 35624 21014 35676 21020
rect 35532 20936 35584 20942
rect 35532 20878 35584 20884
rect 34888 20868 34940 20874
rect 34888 20810 34940 20816
rect 35440 20800 35492 20806
rect 35636 20754 35664 21014
rect 35728 20806 35756 21422
rect 35440 20742 35492 20748
rect 35452 20602 35480 20742
rect 35544 20726 35664 20754
rect 35716 20800 35768 20806
rect 35716 20742 35768 20748
rect 35440 20596 35492 20602
rect 35440 20538 35492 20544
rect 34796 20528 34848 20534
rect 34796 20470 34848 20476
rect 34704 20460 34756 20466
rect 34704 20402 34756 20408
rect 34612 19372 34664 19378
rect 34612 19314 34664 19320
rect 34716 19310 34744 20402
rect 34808 19990 34836 20470
rect 35348 20392 35400 20398
rect 35348 20334 35400 20340
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 34796 19984 34848 19990
rect 34796 19926 34848 19932
rect 34704 19304 34756 19310
rect 34704 19246 34756 19252
rect 34808 19242 34836 19926
rect 35256 19916 35308 19922
rect 35256 19858 35308 19864
rect 34980 19712 35032 19718
rect 34980 19654 35032 19660
rect 35268 19666 35296 19858
rect 35360 19854 35388 20334
rect 35348 19848 35400 19854
rect 35348 19790 35400 19796
rect 35452 19718 35480 20538
rect 35544 20262 35572 20726
rect 35532 20256 35584 20262
rect 35532 20198 35584 20204
rect 35440 19712 35492 19718
rect 34992 19514 35020 19654
rect 35268 19638 35388 19666
rect 35440 19654 35492 19660
rect 34980 19508 35032 19514
rect 34980 19450 35032 19456
rect 35360 19446 35388 19638
rect 35348 19440 35400 19446
rect 35348 19382 35400 19388
rect 34796 19236 34848 19242
rect 34796 19178 34848 19184
rect 34520 18828 34572 18834
rect 34520 18770 34572 18776
rect 34808 18766 34836 19178
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 34980 18828 35032 18834
rect 34980 18770 35032 18776
rect 34796 18760 34848 18766
rect 34796 18702 34848 18708
rect 34992 18426 35020 18770
rect 34980 18420 35032 18426
rect 34980 18362 35032 18368
rect 35360 18290 35388 19382
rect 35544 19174 35572 20198
rect 35532 19168 35584 19174
rect 35532 19110 35584 19116
rect 35348 18284 35400 18290
rect 35348 18226 35400 18232
rect 34060 18216 34112 18222
rect 34060 18158 34112 18164
rect 34336 18216 34388 18222
rect 34336 18158 34388 18164
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 32956 17740 33008 17746
rect 32956 17682 33008 17688
rect 32404 17672 32456 17678
rect 32404 17614 32456 17620
rect 31852 17604 31904 17610
rect 31852 17546 31904 17552
rect 27804 17536 27856 17542
rect 27804 17478 27856 17484
rect 31024 17536 31076 17542
rect 31024 17478 31076 17484
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 25688 16448 25740 16454
rect 25688 16390 25740 16396
rect 25700 16114 25728 16390
rect 25504 16108 25556 16114
rect 25504 16050 25556 16056
rect 25688 16108 25740 16114
rect 25688 16050 25740 16056
rect 26056 16108 26108 16114
rect 26056 16050 26108 16056
rect 23756 15700 23808 15706
rect 23756 15642 23808 15648
rect 25044 15700 25096 15706
rect 25044 15642 25096 15648
rect 23572 15496 23624 15502
rect 25504 15496 25556 15502
rect 23572 15438 23624 15444
rect 25240 15444 25504 15450
rect 25240 15438 25556 15444
rect 25240 15422 25544 15438
rect 23940 15360 23992 15366
rect 23940 15302 23992 15308
rect 23952 15162 23980 15302
rect 23940 15156 23992 15162
rect 23940 15098 23992 15104
rect 23112 15020 23164 15026
rect 23112 14962 23164 14968
rect 23124 14618 23152 14962
rect 23952 14618 23980 15098
rect 25240 14958 25268 15422
rect 25320 15360 25372 15366
rect 25320 15302 25372 15308
rect 25504 15360 25556 15366
rect 25504 15302 25556 15308
rect 25332 15026 25360 15302
rect 25320 15020 25372 15026
rect 25320 14962 25372 14968
rect 24308 14952 24360 14958
rect 24308 14894 24360 14900
rect 25228 14952 25280 14958
rect 25228 14894 25280 14900
rect 25412 14952 25464 14958
rect 25412 14894 25464 14900
rect 23112 14612 23164 14618
rect 23112 14554 23164 14560
rect 23940 14612 23992 14618
rect 23940 14554 23992 14560
rect 24320 14346 24348 14894
rect 25044 14884 25096 14890
rect 25044 14826 25096 14832
rect 25056 14482 25084 14826
rect 25044 14476 25096 14482
rect 25044 14418 25096 14424
rect 24676 14408 24728 14414
rect 24728 14368 24900 14396
rect 24676 14350 24728 14356
rect 24308 14340 24360 14346
rect 24308 14282 24360 14288
rect 24124 14272 24176 14278
rect 24124 14214 24176 14220
rect 22836 14068 22888 14074
rect 22388 14028 22508 14056
rect 22376 13932 22428 13938
rect 22376 13874 22428 13880
rect 22284 13320 22336 13326
rect 22284 13262 22336 13268
rect 22388 13190 22416 13874
rect 22480 13870 22508 14028
rect 22836 14010 22888 14016
rect 24136 13938 24164 14214
rect 24872 14006 24900 14368
rect 25228 14340 25280 14346
rect 25228 14282 25280 14288
rect 24860 14000 24912 14006
rect 24860 13942 24912 13948
rect 24124 13932 24176 13938
rect 24124 13874 24176 13880
rect 24952 13932 25004 13938
rect 24952 13874 25004 13880
rect 25044 13932 25096 13938
rect 25044 13874 25096 13880
rect 22468 13864 22520 13870
rect 22468 13806 22520 13812
rect 23756 13864 23808 13870
rect 23756 13806 23808 13812
rect 24216 13864 24268 13870
rect 24216 13806 24268 13812
rect 23664 13728 23716 13734
rect 23664 13670 23716 13676
rect 22376 13184 22428 13190
rect 22376 13126 22428 13132
rect 23388 13184 23440 13190
rect 23388 13126 23440 13132
rect 22100 12980 22152 12986
rect 22100 12922 22152 12928
rect 22192 12844 22244 12850
rect 22192 12786 22244 12792
rect 22204 12238 22232 12786
rect 23400 12306 23428 13126
rect 23676 12850 23704 13670
rect 23664 12844 23716 12850
rect 23664 12786 23716 12792
rect 23768 12306 23796 13806
rect 24124 13184 24176 13190
rect 24124 13126 24176 13132
rect 24136 12850 24164 13126
rect 24124 12844 24176 12850
rect 24124 12786 24176 12792
rect 24228 12782 24256 13806
rect 24964 13462 24992 13874
rect 24952 13456 25004 13462
rect 24952 13398 25004 13404
rect 25056 13394 25084 13874
rect 25240 13870 25268 14282
rect 25424 14278 25452 14894
rect 25412 14272 25464 14278
rect 25412 14214 25464 14220
rect 25228 13864 25280 13870
rect 25228 13806 25280 13812
rect 25240 13734 25268 13806
rect 25228 13728 25280 13734
rect 25228 13670 25280 13676
rect 25044 13388 25096 13394
rect 25044 13330 25096 13336
rect 24768 13320 24820 13326
rect 24768 13262 24820 13268
rect 24780 12782 24808 13262
rect 24952 13184 25004 13190
rect 24952 13126 25004 13132
rect 24964 12850 24992 13126
rect 24952 12844 25004 12850
rect 24952 12786 25004 12792
rect 24216 12776 24268 12782
rect 24216 12718 24268 12724
rect 24768 12776 24820 12782
rect 24768 12718 24820 12724
rect 23388 12300 23440 12306
rect 23388 12242 23440 12248
rect 23756 12300 23808 12306
rect 23756 12242 23808 12248
rect 22192 12232 22244 12238
rect 22192 12174 22244 12180
rect 23572 12232 23624 12238
rect 23572 12174 23624 12180
rect 21916 11620 21968 11626
rect 21916 11562 21968 11568
rect 21640 11008 21692 11014
rect 21640 10950 21692 10956
rect 21928 10674 21956 11562
rect 22204 11286 22232 12174
rect 22744 12096 22796 12102
rect 22744 12038 22796 12044
rect 22756 11694 22784 12038
rect 23480 11756 23532 11762
rect 23480 11698 23532 11704
rect 22744 11688 22796 11694
rect 22744 11630 22796 11636
rect 22192 11280 22244 11286
rect 22192 11222 22244 11228
rect 23492 11150 23520 11698
rect 23584 11694 23612 12174
rect 24228 11694 24256 12718
rect 24584 12708 24636 12714
rect 24584 12650 24636 12656
rect 24596 12306 24624 12650
rect 24768 12640 24820 12646
rect 24768 12582 24820 12588
rect 24584 12300 24636 12306
rect 24584 12242 24636 12248
rect 23572 11688 23624 11694
rect 23572 11630 23624 11636
rect 24216 11688 24268 11694
rect 24216 11630 24268 11636
rect 23584 11150 23612 11630
rect 24228 11558 24256 11630
rect 24124 11552 24176 11558
rect 24124 11494 24176 11500
rect 24216 11552 24268 11558
rect 24216 11494 24268 11500
rect 23480 11144 23532 11150
rect 23480 11086 23532 11092
rect 23572 11144 23624 11150
rect 23572 11086 23624 11092
rect 23584 10742 23612 11086
rect 23572 10736 23624 10742
rect 23572 10678 23624 10684
rect 21272 10668 21324 10674
rect 21272 10610 21324 10616
rect 21916 10668 21968 10674
rect 21916 10610 21968 10616
rect 20720 10124 20772 10130
rect 20720 10066 20772 10072
rect 20732 9654 20760 10066
rect 20720 9648 20772 9654
rect 20720 9590 20772 9596
rect 20996 9580 21048 9586
rect 20996 9522 21048 9528
rect 21008 9178 21036 9522
rect 21284 9382 21312 10610
rect 21364 10600 21416 10606
rect 21364 10542 21416 10548
rect 21376 9382 21404 10542
rect 21272 9376 21324 9382
rect 21272 9318 21324 9324
rect 21364 9376 21416 9382
rect 21364 9318 21416 9324
rect 20996 9172 21048 9178
rect 20996 9114 21048 9120
rect 20168 9036 20220 9042
rect 20168 8978 20220 8984
rect 19064 8968 19116 8974
rect 19064 8910 19116 8916
rect 21284 8906 21312 9318
rect 21928 9042 21956 10610
rect 22652 10600 22704 10606
rect 22652 10542 22704 10548
rect 22284 10464 22336 10470
rect 22284 10406 22336 10412
rect 22100 9988 22152 9994
rect 22100 9930 22152 9936
rect 22112 9178 22140 9930
rect 22100 9172 22152 9178
rect 22100 9114 22152 9120
rect 21916 9036 21968 9042
rect 21916 8978 21968 8984
rect 22296 8974 22324 10406
rect 22664 10266 22692 10542
rect 22928 10464 22980 10470
rect 22928 10406 22980 10412
rect 22652 10260 22704 10266
rect 22652 10202 22704 10208
rect 22744 9580 22796 9586
rect 22744 9522 22796 9528
rect 22756 9178 22784 9522
rect 22744 9172 22796 9178
rect 22744 9114 22796 9120
rect 22940 8974 22968 10406
rect 24136 10198 24164 11494
rect 24228 10538 24256 11494
rect 24676 11280 24728 11286
rect 24676 11222 24728 11228
rect 24584 11076 24636 11082
rect 24584 11018 24636 11024
rect 24216 10532 24268 10538
rect 24216 10474 24268 10480
rect 24596 10266 24624 11018
rect 24584 10260 24636 10266
rect 24584 10202 24636 10208
rect 24124 10192 24176 10198
rect 24124 10134 24176 10140
rect 24688 10130 24716 11222
rect 24780 11150 24808 12582
rect 25424 12374 25452 14214
rect 25516 14006 25544 15302
rect 25700 15162 25728 16050
rect 26068 15706 26096 16050
rect 26240 15904 26292 15910
rect 26240 15846 26292 15852
rect 26056 15700 26108 15706
rect 26056 15642 26108 15648
rect 25688 15156 25740 15162
rect 25688 15098 25740 15104
rect 25700 14482 25728 15098
rect 26068 15026 26096 15642
rect 26056 15020 26108 15026
rect 26056 14962 26108 14968
rect 25964 14816 26016 14822
rect 25964 14758 26016 14764
rect 25688 14476 25740 14482
rect 25688 14418 25740 14424
rect 25504 14000 25556 14006
rect 25504 13942 25556 13948
rect 25516 13190 25544 13942
rect 25976 13734 26004 14758
rect 26252 14414 26280 15846
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 26240 14408 26292 14414
rect 26240 14350 26292 14356
rect 26516 14068 26568 14074
rect 26516 14010 26568 14016
rect 26056 14000 26108 14006
rect 26056 13942 26108 13948
rect 25964 13728 26016 13734
rect 25964 13670 26016 13676
rect 25596 13456 25648 13462
rect 25596 13398 25648 13404
rect 25504 13184 25556 13190
rect 25504 13126 25556 13132
rect 25412 12368 25464 12374
rect 25412 12310 25464 12316
rect 25320 11552 25372 11558
rect 25320 11494 25372 11500
rect 24768 11144 24820 11150
rect 24768 11086 24820 11092
rect 24676 10124 24728 10130
rect 24676 10066 24728 10072
rect 25332 10062 25360 11494
rect 25412 11076 25464 11082
rect 25412 11018 25464 11024
rect 25424 10266 25452 11018
rect 25608 11014 25636 13398
rect 25688 13252 25740 13258
rect 25688 13194 25740 13200
rect 25700 12434 25728 13194
rect 25780 13184 25832 13190
rect 25780 13126 25832 13132
rect 25792 12782 25820 13126
rect 25780 12776 25832 12782
rect 25780 12718 25832 12724
rect 25792 12594 25820 12718
rect 25792 12566 26004 12594
rect 25700 12406 25912 12434
rect 25884 12238 25912 12406
rect 25872 12232 25924 12238
rect 25700 12192 25872 12220
rect 25700 11218 25728 12192
rect 25872 12174 25924 12180
rect 25976 11694 26004 12566
rect 26068 11762 26096 13942
rect 26148 13728 26200 13734
rect 26148 13670 26200 13676
rect 26424 13728 26476 13734
rect 26424 13670 26476 13676
rect 26160 13546 26188 13670
rect 26160 13518 26372 13546
rect 26148 13456 26200 13462
rect 26148 13398 26200 13404
rect 26160 13258 26188 13398
rect 26344 13394 26372 13518
rect 26332 13388 26384 13394
rect 26332 13330 26384 13336
rect 26148 13252 26200 13258
rect 26148 13194 26200 13200
rect 26332 13252 26384 13258
rect 26332 13194 26384 13200
rect 26344 12986 26372 13194
rect 26332 12980 26384 12986
rect 26332 12922 26384 12928
rect 26240 12912 26292 12918
rect 26160 12860 26240 12866
rect 26160 12854 26292 12860
rect 26160 12838 26280 12854
rect 26436 12850 26464 13670
rect 26424 12844 26476 12850
rect 26160 12186 26188 12838
rect 26424 12786 26476 12792
rect 26528 12782 26556 14010
rect 26792 13796 26844 13802
rect 26792 13738 26844 13744
rect 27620 13796 27672 13802
rect 27620 13738 27672 13744
rect 26804 12782 26832 13738
rect 26976 13320 27028 13326
rect 26976 13262 27028 13268
rect 26988 12850 27016 13262
rect 27160 13252 27212 13258
rect 27160 13194 27212 13200
rect 27172 12850 27200 13194
rect 27632 13190 27660 13738
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 27620 13184 27672 13190
rect 27620 13126 27672 13132
rect 27632 12918 27660 13126
rect 27620 12912 27672 12918
rect 27620 12854 27672 12860
rect 26976 12844 27028 12850
rect 26976 12786 27028 12792
rect 27160 12844 27212 12850
rect 27160 12786 27212 12792
rect 28172 12844 28224 12850
rect 28172 12786 28224 12792
rect 26516 12776 26568 12782
rect 26516 12718 26568 12724
rect 26792 12776 26844 12782
rect 26792 12718 26844 12724
rect 26240 12708 26292 12714
rect 26240 12650 26292 12656
rect 26252 12374 26280 12650
rect 26240 12368 26292 12374
rect 26240 12310 26292 12316
rect 26424 12232 26476 12238
rect 26160 12180 26424 12186
rect 26528 12220 26556 12718
rect 26608 12232 26660 12238
rect 26528 12192 26608 12220
rect 26160 12174 26476 12180
rect 26608 12174 26660 12180
rect 26160 12158 26464 12174
rect 26056 11756 26108 11762
rect 26056 11698 26108 11704
rect 25964 11688 26016 11694
rect 25964 11630 26016 11636
rect 25688 11212 25740 11218
rect 25688 11154 25740 11160
rect 25596 11008 25648 11014
rect 25596 10950 25648 10956
rect 25412 10260 25464 10266
rect 25412 10202 25464 10208
rect 25608 10130 25636 10950
rect 25700 10674 25728 11154
rect 25976 11082 26004 11630
rect 26160 11558 26188 12158
rect 26424 11756 26476 11762
rect 26424 11698 26476 11704
rect 26240 11688 26292 11694
rect 26240 11630 26292 11636
rect 26148 11552 26200 11558
rect 26148 11494 26200 11500
rect 26252 11218 26280 11630
rect 26332 11552 26384 11558
rect 26332 11494 26384 11500
rect 26240 11212 26292 11218
rect 26240 11154 26292 11160
rect 25964 11076 26016 11082
rect 25964 11018 26016 11024
rect 26148 11008 26200 11014
rect 26148 10950 26200 10956
rect 25688 10668 25740 10674
rect 25688 10610 25740 10616
rect 25596 10124 25648 10130
rect 25596 10066 25648 10072
rect 25700 10062 25728 10610
rect 26160 10538 26188 10950
rect 26344 10674 26372 11494
rect 26436 11286 26464 11698
rect 26804 11626 26832 12718
rect 27068 12232 27120 12238
rect 27068 12174 27120 12180
rect 27080 11762 27108 12174
rect 27172 11898 27200 12786
rect 28184 12442 28212 12786
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 27620 12436 27672 12442
rect 27620 12378 27672 12384
rect 28172 12436 28224 12442
rect 28172 12378 28224 12384
rect 27160 11892 27212 11898
rect 27160 11834 27212 11840
rect 27632 11762 27660 12378
rect 27068 11756 27120 11762
rect 27068 11698 27120 11704
rect 27620 11756 27672 11762
rect 27620 11698 27672 11704
rect 26792 11620 26844 11626
rect 26792 11562 26844 11568
rect 26424 11280 26476 11286
rect 26424 11222 26476 11228
rect 26516 11212 26568 11218
rect 26516 11154 26568 11160
rect 26608 11212 26660 11218
rect 26608 11154 26660 11160
rect 26332 10668 26384 10674
rect 26332 10610 26384 10616
rect 26528 10606 26556 11154
rect 26516 10600 26568 10606
rect 26516 10542 26568 10548
rect 26148 10532 26200 10538
rect 26148 10474 26200 10480
rect 25320 10056 25372 10062
rect 25320 9998 25372 10004
rect 25688 10056 25740 10062
rect 25688 9998 25740 10004
rect 22284 8968 22336 8974
rect 22284 8910 22336 8916
rect 22928 8968 22980 8974
rect 22928 8910 22980 8916
rect 18052 8900 18104 8906
rect 18052 8842 18104 8848
rect 21272 8900 21324 8906
rect 21272 8842 21324 8848
rect 18604 8832 18656 8838
rect 18604 8774 18656 8780
rect 17592 8492 17644 8498
rect 17592 8434 17644 8440
rect 17316 8288 17368 8294
rect 17316 8230 17368 8236
rect 17224 8084 17276 8090
rect 17224 8026 17276 8032
rect 16580 7948 16632 7954
rect 16580 7890 16632 7896
rect 11520 7880 11572 7886
rect 11520 7822 11572 7828
rect 12532 7880 12584 7886
rect 12532 7822 12584 7828
rect 17236 7410 17264 8026
rect 17328 7886 17356 8230
rect 17316 7880 17368 7886
rect 17316 7822 17368 7828
rect 17604 7546 17632 8434
rect 18616 8090 18644 8774
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 18604 8084 18656 8090
rect 18604 8026 18656 8032
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 17592 7540 17644 7546
rect 17592 7482 17644 7488
rect 17224 7404 17276 7410
rect 17224 7346 17276 7352
rect 17408 7404 17460 7410
rect 17408 7346 17460 7352
rect 11336 6792 11388 6798
rect 11336 6734 11388 6740
rect 9220 2644 9272 2650
rect 9220 2586 9272 2592
rect 11244 2644 11296 2650
rect 11244 2586 11296 2592
rect 17420 2514 17448 7346
rect 26620 6914 26648 11154
rect 26804 11150 26832 11562
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 26792 11144 26844 11150
rect 26792 11086 26844 11092
rect 35820 10470 35848 37198
rect 38200 34604 38252 34610
rect 38200 34546 38252 34552
rect 38016 34400 38068 34406
rect 38016 34342 38068 34348
rect 38028 34105 38056 34342
rect 38014 34096 38070 34105
rect 38014 34031 38070 34040
rect 36084 31952 36136 31958
rect 36084 31894 36136 31900
rect 35992 31204 36044 31210
rect 35992 31146 36044 31152
rect 36004 30802 36032 31146
rect 35992 30796 36044 30802
rect 35992 30738 36044 30744
rect 35900 30728 35952 30734
rect 35900 30670 35952 30676
rect 35912 30054 35940 30670
rect 35900 30048 35952 30054
rect 35900 29990 35952 29996
rect 35900 28960 35952 28966
rect 35900 28902 35952 28908
rect 35912 28558 35940 28902
rect 35900 28552 35952 28558
rect 35900 28494 35952 28500
rect 35912 28082 35940 28494
rect 35992 28484 36044 28490
rect 35992 28426 36044 28432
rect 36004 28082 36032 28426
rect 35900 28076 35952 28082
rect 35900 28018 35952 28024
rect 35992 28076 36044 28082
rect 35992 28018 36044 28024
rect 36004 27538 36032 28018
rect 36096 27577 36124 31894
rect 36176 30592 36228 30598
rect 36176 30534 36228 30540
rect 37188 30592 37240 30598
rect 37188 30534 37240 30540
rect 36188 30190 36216 30534
rect 36268 30252 36320 30258
rect 36268 30194 36320 30200
rect 36176 30184 36228 30190
rect 36176 30126 36228 30132
rect 36188 29646 36216 30126
rect 36280 29782 36308 30194
rect 36544 30048 36596 30054
rect 36544 29990 36596 29996
rect 36268 29776 36320 29782
rect 36268 29718 36320 29724
rect 36176 29640 36228 29646
rect 36176 29582 36228 29588
rect 36280 29578 36308 29718
rect 36268 29572 36320 29578
rect 36268 29514 36320 29520
rect 36556 29238 36584 29990
rect 36544 29232 36596 29238
rect 36544 29174 36596 29180
rect 36556 28558 36584 29174
rect 36636 29164 36688 29170
rect 36636 29106 36688 29112
rect 36544 28552 36596 28558
rect 36544 28494 36596 28500
rect 36544 28416 36596 28422
rect 36544 28358 36596 28364
rect 36556 28082 36584 28358
rect 36544 28076 36596 28082
rect 36544 28018 36596 28024
rect 36648 28014 36676 29106
rect 36636 28008 36688 28014
rect 36636 27950 36688 27956
rect 36636 27872 36688 27878
rect 36636 27814 36688 27820
rect 36082 27568 36138 27577
rect 35992 27532 36044 27538
rect 36358 27568 36414 27577
rect 36082 27503 36138 27512
rect 36176 27532 36228 27538
rect 35992 27474 36044 27480
rect 36358 27503 36414 27512
rect 36176 27474 36228 27480
rect 36084 27328 36136 27334
rect 36084 27270 36136 27276
rect 35900 26988 35952 26994
rect 35900 26930 35952 26936
rect 35912 26625 35940 26930
rect 35898 26616 35954 26625
rect 35898 26551 35900 26560
rect 35952 26551 35954 26560
rect 35900 26522 35952 26528
rect 36096 26466 36124 27270
rect 36188 26586 36216 27474
rect 36372 27470 36400 27503
rect 36360 27464 36412 27470
rect 36360 27406 36412 27412
rect 36450 27024 36506 27033
rect 36450 26959 36452 26968
rect 36504 26959 36506 26968
rect 36544 26988 36596 26994
rect 36452 26930 36504 26936
rect 36544 26930 36596 26936
rect 36452 26784 36504 26790
rect 36452 26726 36504 26732
rect 36176 26580 36228 26586
rect 36176 26522 36228 26528
rect 36096 26438 36216 26466
rect 36188 25906 36216 26438
rect 36464 26382 36492 26726
rect 36452 26376 36504 26382
rect 36452 26318 36504 26324
rect 36556 26246 36584 26930
rect 36544 26240 36596 26246
rect 36544 26182 36596 26188
rect 35992 25900 36044 25906
rect 35992 25842 36044 25848
rect 36176 25900 36228 25906
rect 36176 25842 36228 25848
rect 35900 25696 35952 25702
rect 35900 25638 35952 25644
rect 35912 24886 35940 25638
rect 36004 25158 36032 25842
rect 36188 25498 36216 25842
rect 36176 25492 36228 25498
rect 36176 25434 36228 25440
rect 35992 25152 36044 25158
rect 35992 25094 36044 25100
rect 36176 25152 36228 25158
rect 36176 25094 36228 25100
rect 35900 24880 35952 24886
rect 35900 24822 35952 24828
rect 36004 24818 36032 25094
rect 35992 24812 36044 24818
rect 35992 24754 36044 24760
rect 36188 24750 36216 25094
rect 36176 24744 36228 24750
rect 36176 24686 36228 24692
rect 36268 24608 36320 24614
rect 36268 24550 36320 24556
rect 35900 23792 35952 23798
rect 35900 23734 35952 23740
rect 35912 22982 35940 23734
rect 35900 22976 35952 22982
rect 35900 22918 35952 22924
rect 36084 22976 36136 22982
rect 36084 22918 36136 22924
rect 36096 22642 36124 22918
rect 36280 22642 36308 24550
rect 36648 23798 36676 27814
rect 36728 27532 36780 27538
rect 36728 27474 36780 27480
rect 36740 26858 36768 27474
rect 37200 26994 37228 30534
rect 37924 30252 37976 30258
rect 37924 30194 37976 30200
rect 37372 30184 37424 30190
rect 37372 30126 37424 30132
rect 37384 29850 37412 30126
rect 37832 30116 37884 30122
rect 37832 30058 37884 30064
rect 37372 29844 37424 29850
rect 37372 29786 37424 29792
rect 37280 29096 37332 29102
rect 37280 29038 37332 29044
rect 37464 29096 37516 29102
rect 37464 29038 37516 29044
rect 37292 28762 37320 29038
rect 37280 28756 37332 28762
rect 37280 28698 37332 28704
rect 37280 28552 37332 28558
rect 37280 28494 37332 28500
rect 37292 28082 37320 28494
rect 37476 28490 37504 29038
rect 37648 28756 37700 28762
rect 37648 28698 37700 28704
rect 37464 28484 37516 28490
rect 37464 28426 37516 28432
rect 37372 28416 37424 28422
rect 37372 28358 37424 28364
rect 37280 28076 37332 28082
rect 37280 28018 37332 28024
rect 37280 27328 37332 27334
rect 37280 27270 37332 27276
rect 37188 26988 37240 26994
rect 37188 26930 37240 26936
rect 36728 26852 36780 26858
rect 36728 26794 36780 26800
rect 36740 26042 36768 26794
rect 36728 26036 36780 26042
rect 36728 25978 36780 25984
rect 36728 24812 36780 24818
rect 36728 24754 36780 24760
rect 36740 24410 36768 24754
rect 37188 24744 37240 24750
rect 37188 24686 37240 24692
rect 36728 24404 36780 24410
rect 36728 24346 36780 24352
rect 37096 24200 37148 24206
rect 37096 24142 37148 24148
rect 36636 23792 36688 23798
rect 36636 23734 36688 23740
rect 36728 23520 36780 23526
rect 36728 23462 36780 23468
rect 36740 23322 36768 23462
rect 37108 23322 37136 24142
rect 37200 23730 37228 24686
rect 37292 24274 37320 27270
rect 37384 26926 37412 28358
rect 37476 28082 37504 28426
rect 37660 28218 37688 28698
rect 37648 28212 37700 28218
rect 37648 28154 37700 28160
rect 37464 28076 37516 28082
rect 37464 28018 37516 28024
rect 37476 27606 37504 28018
rect 37740 27872 37792 27878
rect 37740 27814 37792 27820
rect 37464 27600 37516 27606
rect 37464 27542 37516 27548
rect 37752 27470 37780 27814
rect 37740 27464 37792 27470
rect 37740 27406 37792 27412
rect 37372 26920 37424 26926
rect 37372 26862 37424 26868
rect 37740 26784 37792 26790
rect 37740 26726 37792 26732
rect 37556 26512 37608 26518
rect 37556 26454 37608 26460
rect 37372 26308 37424 26314
rect 37372 26250 37424 26256
rect 37280 24268 37332 24274
rect 37280 24210 37332 24216
rect 37292 24138 37320 24210
rect 37280 24132 37332 24138
rect 37280 24074 37332 24080
rect 37188 23724 37240 23730
rect 37188 23666 37240 23672
rect 36728 23316 36780 23322
rect 36728 23258 36780 23264
rect 37096 23316 37148 23322
rect 37096 23258 37148 23264
rect 36636 23112 36688 23118
rect 36636 23054 36688 23060
rect 36084 22636 36136 22642
rect 36084 22578 36136 22584
rect 36268 22636 36320 22642
rect 36268 22578 36320 22584
rect 36648 22506 36676 23054
rect 35900 22500 35952 22506
rect 35900 22442 35952 22448
rect 36636 22500 36688 22506
rect 36636 22442 36688 22448
rect 35912 21554 35940 22442
rect 36740 22438 36768 23258
rect 36728 22432 36780 22438
rect 36728 22374 36780 22380
rect 37384 22030 37412 26250
rect 37464 25900 37516 25906
rect 37464 25842 37516 25848
rect 37476 24954 37504 25842
rect 37568 25838 37596 26454
rect 37752 26382 37780 26726
rect 37740 26376 37792 26382
rect 37740 26318 37792 26324
rect 37556 25832 37608 25838
rect 37556 25774 37608 25780
rect 37556 25696 37608 25702
rect 37556 25638 37608 25644
rect 37568 25362 37596 25638
rect 37556 25356 37608 25362
rect 37556 25298 37608 25304
rect 37844 25294 37872 30058
rect 37936 29306 37964 30194
rect 37924 29300 37976 29306
rect 37924 29242 37976 29248
rect 37924 29028 37976 29034
rect 37924 28970 37976 28976
rect 37936 28490 37964 28970
rect 37924 28484 37976 28490
rect 37924 28426 37976 28432
rect 37936 28082 37964 28426
rect 38108 28416 38160 28422
rect 38108 28358 38160 28364
rect 37924 28076 37976 28082
rect 37924 28018 37976 28024
rect 38120 27470 38148 28358
rect 38108 27464 38160 27470
rect 38108 27406 38160 27412
rect 37832 25288 37884 25294
rect 37832 25230 37884 25236
rect 37556 25152 37608 25158
rect 37556 25094 37608 25100
rect 37464 24948 37516 24954
rect 37464 24890 37516 24896
rect 37372 22024 37424 22030
rect 37372 21966 37424 21972
rect 35900 21548 35952 21554
rect 35900 21490 35952 21496
rect 36084 21548 36136 21554
rect 36084 21490 36136 21496
rect 35912 21078 35940 21490
rect 35992 21412 36044 21418
rect 35992 21354 36044 21360
rect 36004 21078 36032 21354
rect 35900 21072 35952 21078
rect 35900 21014 35952 21020
rect 35992 21072 36044 21078
rect 35992 21014 36044 21020
rect 35900 20936 35952 20942
rect 35900 20878 35952 20884
rect 35912 20806 35940 20878
rect 35900 20800 35952 20806
rect 35900 20742 35952 20748
rect 36004 20398 36032 21014
rect 36096 20942 36124 21490
rect 37568 21486 37596 25094
rect 37740 24812 37792 24818
rect 37660 24772 37740 24800
rect 37660 23322 37688 24772
rect 37740 24754 37792 24760
rect 37740 24064 37792 24070
rect 37740 24006 37792 24012
rect 37752 23662 37780 24006
rect 37740 23656 37792 23662
rect 37740 23598 37792 23604
rect 37648 23316 37700 23322
rect 37648 23258 37700 23264
rect 37752 23118 37780 23598
rect 37832 23520 37884 23526
rect 37832 23462 37884 23468
rect 37740 23112 37792 23118
rect 37740 23054 37792 23060
rect 37740 22024 37792 22030
rect 37740 21966 37792 21972
rect 37752 21690 37780 21966
rect 37740 21684 37792 21690
rect 37740 21626 37792 21632
rect 37648 21548 37700 21554
rect 37648 21490 37700 21496
rect 37556 21480 37608 21486
rect 37556 21422 37608 21428
rect 37660 21146 37688 21490
rect 37648 21140 37700 21146
rect 37648 21082 37700 21088
rect 37844 21078 37872 23462
rect 38108 21888 38160 21894
rect 38108 21830 38160 21836
rect 38120 21593 38148 21830
rect 38106 21584 38162 21593
rect 38106 21519 38162 21528
rect 37832 21072 37884 21078
rect 37832 21014 37884 21020
rect 36084 20936 36136 20942
rect 36084 20878 36136 20884
rect 36176 20460 36228 20466
rect 36176 20402 36228 20408
rect 35992 20392 36044 20398
rect 35992 20334 36044 20340
rect 36188 20058 36216 20402
rect 36176 20052 36228 20058
rect 36176 19994 36228 20000
rect 37740 14272 37792 14278
rect 37740 14214 37792 14220
rect 35808 10464 35860 10470
rect 35808 10406 35860 10412
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 26528 6886 26648 6914
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 17408 2508 17460 2514
rect 17408 2450 17460 2456
rect 26528 2446 26556 6886
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 37752 2446 37780 14214
rect 37832 12844 37884 12850
rect 37832 12786 37884 12792
rect 37844 12170 37872 12786
rect 38212 12714 38240 34546
rect 38200 12708 38252 12714
rect 38200 12650 38252 12656
rect 38016 12640 38068 12646
rect 38016 12582 38068 12588
rect 38028 12345 38056 12582
rect 38014 12336 38070 12345
rect 38014 12271 38070 12280
rect 37832 12164 37884 12170
rect 37832 12106 37884 12112
rect 20 2440 72 2446
rect 20 2382 72 2388
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 26516 2440 26568 2446
rect 26516 2382 26568 2388
rect 30932 2440 30984 2446
rect 30932 2382 30984 2388
rect 37740 2440 37792 2446
rect 37740 2382 37792 2388
rect 32 800 60 2382
rect 10336 800 10364 2382
rect 20628 2304 20680 2310
rect 20628 2246 20680 2252
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 20640 800 20668 2246
rect 30944 800 30972 2382
rect 38016 2304 38068 2310
rect 38016 2246 38068 2252
rect 38028 1465 38056 2246
rect 38014 1456 38070 1465
rect 38014 1391 38070 1400
rect 18 0 74 800
rect 10322 0 10378 800
rect 20626 0 20682 800
rect 30930 0 30986 800
<< via2 >>
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 1398 21800 1454 21856
rect 1582 32716 1584 32736
rect 1584 32716 1636 32736
rect 1636 32716 1638 32736
rect 1582 32680 1638 32716
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 11610 24148 11612 24168
rect 11612 24148 11664 24168
rect 11664 24148 11666 24168
rect 11610 24112 11666 24148
rect 9678 19352 9734 19408
rect 10414 19488 10470 19544
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 10598 19388 10600 19408
rect 10600 19388 10652 19408
rect 10652 19388 10654 19408
rect 10598 19352 10654 19388
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 9954 12416 10010 12472
rect 1582 10956 1584 10976
rect 1584 10956 1636 10976
rect 1636 10956 1638 10976
rect 1582 10920 1638 10956
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 12346 19488 12402 19544
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19522 30676 19524 30696
rect 19524 30676 19576 30696
rect 19576 30676 19578 30696
rect 19522 30640 19578 30676
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 20442 30640 20498 30696
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 15014 24132 15070 24168
rect 15014 24112 15016 24132
rect 15016 24112 15068 24132
rect 15068 24112 15070 24132
rect 15382 21564 15384 21584
rect 15384 21564 15436 21584
rect 15436 21564 15438 21584
rect 15382 21528 15438 21564
rect 15842 21936 15898 21992
rect 15290 18672 15346 18728
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 14738 13268 14740 13288
rect 14740 13268 14792 13288
rect 14792 13268 14794 13288
rect 14738 13232 14794 13268
rect 15750 13268 15752 13288
rect 15752 13268 15804 13288
rect 15804 13268 15806 13288
rect 15750 13232 15806 13268
rect 18694 26968 18750 27024
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19522 26868 19524 26888
rect 19524 26868 19576 26888
rect 19576 26868 19578 26888
rect 19522 26832 19578 26868
rect 20166 27412 20168 27432
rect 20168 27412 20220 27432
rect 20220 27412 20222 27432
rect 20166 27376 20222 27412
rect 20718 27376 20774 27432
rect 20442 27104 20498 27160
rect 20166 26696 20222 26752
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 18326 21528 18382 21584
rect 18602 21548 18658 21584
rect 18602 21528 18604 21548
rect 18604 21528 18656 21548
rect 18656 21528 18658 21548
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 18418 18672 18474 18728
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 20534 24812 20590 24848
rect 20534 24792 20536 24812
rect 20536 24792 20588 24812
rect 20588 24792 20590 24812
rect 20442 24268 20498 24304
rect 20442 24248 20444 24268
rect 20444 24248 20496 24268
rect 20496 24248 20498 24268
rect 20442 24132 20498 24168
rect 20442 24112 20444 24132
rect 20444 24112 20496 24132
rect 20496 24112 20498 24132
rect 21178 23976 21234 24032
rect 21086 23568 21142 23624
rect 21546 23296 21602 23352
rect 21822 24556 21824 24576
rect 21824 24556 21876 24576
rect 21876 24556 21878 24576
rect 21822 24520 21878 24556
rect 20442 21936 20498 21992
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19798 19388 19800 19408
rect 19800 19388 19852 19408
rect 19852 19388 19854 19408
rect 19798 19352 19854 19388
rect 19798 19252 19800 19272
rect 19800 19252 19852 19272
rect 19852 19252 19854 19272
rect 19798 19216 19854 19252
rect 19706 18808 19762 18864
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 17222 12436 17278 12472
rect 17222 12416 17224 12436
rect 17224 12416 17276 12436
rect 17276 12416 17278 12436
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 20166 19488 20222 19544
rect 20350 19508 20406 19544
rect 20350 19488 20352 19508
rect 20352 19488 20404 19508
rect 20404 19488 20406 19508
rect 22834 28872 22890 28928
rect 22374 26988 22430 27024
rect 22374 26968 22376 26988
rect 22376 26968 22428 26988
rect 22428 26968 22430 26988
rect 22190 24520 22246 24576
rect 22098 23840 22154 23896
rect 22466 23604 22468 23624
rect 22468 23604 22520 23624
rect 22520 23604 22522 23624
rect 22466 23568 22522 23604
rect 22742 24556 22744 24576
rect 22744 24556 22796 24576
rect 22796 24556 22798 24576
rect 22742 24520 22798 24556
rect 22742 23840 22798 23896
rect 20534 19236 20590 19272
rect 20534 19216 20536 19236
rect 20536 19216 20588 19236
rect 20588 19216 20590 19236
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 22006 21528 22062 21584
rect 21822 14340 21878 14376
rect 21822 14320 21824 14340
rect 21824 14320 21876 14340
rect 21876 14320 21878 14340
rect 23018 29844 23074 29880
rect 23018 29824 23020 29844
rect 23020 29824 23072 29844
rect 23072 29824 23074 29844
rect 22742 14356 22744 14376
rect 22744 14356 22796 14376
rect 22796 14356 22798 14376
rect 22742 14320 22798 14356
rect 23662 20052 23718 20088
rect 23662 20032 23664 20052
rect 23664 20032 23716 20052
rect 23716 20032 23718 20052
rect 24214 24248 24270 24304
rect 24398 24248 24454 24304
rect 24306 24012 24308 24032
rect 24308 24012 24360 24032
rect 24360 24012 24362 24032
rect 24306 23976 24362 24012
rect 24306 21548 24362 21584
rect 24306 21528 24308 21548
rect 24308 21528 24360 21548
rect 24360 21528 24362 21548
rect 23478 19760 23534 19816
rect 23662 19352 23718 19408
rect 24950 24112 25006 24168
rect 24306 18828 24362 18864
rect 24306 18808 24308 18828
rect 24308 18808 24360 18828
rect 24360 18808 24362 18828
rect 25410 27104 25466 27160
rect 25318 26988 25374 27024
rect 25318 26968 25320 26988
rect 25320 26968 25372 26988
rect 25372 26968 25374 26988
rect 25686 27104 25742 27160
rect 25870 25764 25926 25800
rect 25870 25744 25872 25764
rect 25872 25744 25924 25764
rect 25924 25744 25926 25764
rect 26238 24812 26294 24848
rect 26238 24792 26240 24812
rect 26240 24792 26292 24812
rect 26292 24792 26294 24812
rect 25870 21664 25926 21720
rect 25778 19236 25834 19272
rect 25778 19216 25780 19236
rect 25780 19216 25832 19236
rect 25832 19216 25834 19236
rect 26422 24520 26478 24576
rect 26054 20032 26110 20088
rect 27066 26424 27122 26480
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 27434 27820 27436 27840
rect 27436 27820 27488 27840
rect 27488 27820 27490 27840
rect 27434 27784 27490 27820
rect 27434 26968 27490 27024
rect 28262 29824 28318 29880
rect 28078 28464 28134 28520
rect 27894 27668 27950 27704
rect 27894 27648 27896 27668
rect 27896 27648 27948 27668
rect 27948 27648 27950 27668
rect 28078 27548 28080 27568
rect 28080 27548 28132 27568
rect 28132 27548 28134 27568
rect 28078 27512 28134 27548
rect 28078 26832 28134 26888
rect 27986 24284 27988 24304
rect 27988 24284 28040 24304
rect 28040 24284 28042 24304
rect 27986 24248 28042 24284
rect 28446 28872 28502 28928
rect 28446 27820 28448 27840
rect 28448 27820 28500 27840
rect 28500 27820 28502 27840
rect 28446 27784 28502 27820
rect 28446 27668 28502 27704
rect 28446 27648 28448 27668
rect 28448 27648 28500 27668
rect 28500 27648 28502 27668
rect 28262 25744 28318 25800
rect 28170 23840 28226 23896
rect 27434 20576 27490 20632
rect 27342 19624 27398 19680
rect 27986 20576 28042 20632
rect 27986 19760 28042 19816
rect 29090 29180 29092 29200
rect 29092 29180 29144 29200
rect 29144 29180 29146 29200
rect 29090 29144 29146 29180
rect 28906 28872 28962 28928
rect 29182 28192 29238 28248
rect 28998 27820 29000 27840
rect 29000 27820 29052 27840
rect 29052 27820 29054 27840
rect 28998 27784 29054 27820
rect 28814 26696 28870 26752
rect 29182 27920 29238 27976
rect 29366 27920 29422 27976
rect 29642 27820 29644 27840
rect 29644 27820 29696 27840
rect 29696 27820 29698 27840
rect 29642 27784 29698 27820
rect 29642 27648 29698 27704
rect 28906 19624 28962 19680
rect 28722 19236 28778 19272
rect 28722 19216 28724 19236
rect 28724 19216 28776 19236
rect 28776 19216 28778 19236
rect 29642 26696 29698 26752
rect 29366 23296 29422 23352
rect 30562 31728 30618 31784
rect 30010 27376 30066 27432
rect 30102 26560 30158 26616
rect 30010 26324 30012 26344
rect 30012 26324 30064 26344
rect 30064 26324 30066 26344
rect 30010 26288 30066 26324
rect 30746 31864 30802 31920
rect 30746 31456 30802 31512
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 30930 32000 30986 32056
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 31482 32000 31538 32056
rect 30930 28600 30986 28656
rect 31114 28328 31170 28384
rect 30838 27784 30894 27840
rect 30930 26152 30986 26208
rect 30746 24928 30802 24984
rect 30930 25200 30986 25256
rect 30746 21664 30802 21720
rect 30562 21528 30618 21584
rect 29642 19388 29644 19408
rect 29644 19388 29696 19408
rect 29696 19388 29698 19408
rect 29642 19352 29698 19388
rect 30378 19352 30434 19408
rect 31482 27512 31538 27568
rect 31482 27276 31484 27296
rect 31484 27276 31536 27296
rect 31536 27276 31538 27296
rect 31482 27240 31538 27276
rect 31390 26968 31446 27024
rect 32034 28500 32036 28520
rect 32036 28500 32088 28520
rect 32088 28500 32090 28520
rect 32034 28464 32090 28500
rect 31850 28092 31852 28112
rect 31852 28092 31904 28112
rect 31904 28092 31906 28112
rect 31850 28056 31906 28092
rect 32126 28192 32182 28248
rect 31942 27668 31998 27704
rect 31942 27648 31944 27668
rect 31944 27648 31996 27668
rect 31996 27648 31998 27668
rect 31850 27548 31852 27568
rect 31852 27548 31904 27568
rect 31904 27548 31906 27568
rect 31850 27512 31906 27548
rect 31850 27240 31906 27296
rect 32034 26968 32090 27024
rect 32678 28192 32734 28248
rect 32218 27648 32274 27704
rect 32586 27784 32642 27840
rect 32402 27376 32458 27432
rect 32494 26832 32550 26888
rect 32954 28328 33010 28384
rect 32862 26560 32918 26616
rect 33414 28328 33470 28384
rect 33230 28056 33286 28112
rect 33322 27240 33378 27296
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 33966 28600 34022 28656
rect 33690 27920 33746 27976
rect 33598 26424 33654 26480
rect 33782 26696 33838 26752
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34150 29144 34206 29200
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34794 27920 34850 27976
rect 34058 26288 34114 26344
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 35346 26560 35402 26616
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 35714 27104 35770 27160
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34518 23160 34574 23216
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 38014 34040 38070 34096
rect 36082 27512 36138 27568
rect 36358 27512 36414 27568
rect 35898 26580 35954 26616
rect 35898 26560 35900 26580
rect 35900 26560 35952 26580
rect 35952 26560 35954 26580
rect 36450 26988 36506 27024
rect 36450 26968 36452 26988
rect 36452 26968 36504 26988
rect 36504 26968 36506 26988
rect 38106 21528 38162 21584
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 38014 12280 38070 12336
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 38014 1400 38070 1456
<< metal3 >>
rect 4208 37568 4528 37569
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 35327 35248 35328
rect 19568 34848 19888 34849
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 4208 34304 4528 34305
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 38009 34098 38075 34101
rect 39200 34098 40000 34128
rect 38009 34096 40000 34098
rect 38009 34040 38014 34096
rect 38070 34040 40000 34096
rect 38009 34038 40000 34040
rect 38009 34035 38075 34038
rect 39200 34008 40000 34038
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 0 32738 800 32768
rect 1577 32738 1643 32741
rect 0 32736 1643 32738
rect 0 32680 1582 32736
rect 1638 32680 1643 32736
rect 0 32678 1643 32680
rect 0 32648 800 32678
rect 1577 32675 1643 32678
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 32607 19888 32608
rect 4208 32128 4528 32129
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 30925 32058 30991 32061
rect 31477 32058 31543 32061
rect 30925 32056 31543 32058
rect 30925 32000 30930 32056
rect 30986 32000 31482 32056
rect 31538 32000 31543 32056
rect 30925 31998 31543 32000
rect 30925 31995 30991 31998
rect 31477 31995 31543 31998
rect 30741 31924 30807 31925
rect 30741 31920 30788 31924
rect 30852 31922 30858 31924
rect 30741 31864 30746 31920
rect 30741 31860 30788 31864
rect 30852 31862 30898 31922
rect 30852 31860 30858 31862
rect 30741 31859 30807 31860
rect 30557 31786 30623 31789
rect 30557 31784 30850 31786
rect 30557 31728 30562 31784
rect 30618 31728 30850 31784
rect 30557 31726 30850 31728
rect 30557 31723 30623 31726
rect 30790 31650 30850 31726
rect 30966 31650 30972 31652
rect 30790 31590 30972 31650
rect 30966 31588 30972 31590
rect 31036 31588 31042 31652
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 30741 31516 30807 31517
rect 30741 31514 30788 31516
rect 30696 31512 30788 31514
rect 30696 31456 30746 31512
rect 30696 31454 30788 31456
rect 30741 31452 30788 31454
rect 30852 31452 30858 31516
rect 30741 31451 30807 31452
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 19517 30698 19583 30701
rect 20437 30698 20503 30701
rect 19517 30696 20503 30698
rect 19517 30640 19522 30696
rect 19578 30640 20442 30696
rect 20498 30640 20503 30696
rect 19517 30638 20503 30640
rect 19517 30635 19583 30638
rect 20437 30635 20503 30638
rect 19568 30496 19888 30497
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 29887 35248 29888
rect 23013 29882 23079 29885
rect 28257 29882 28323 29885
rect 23013 29880 28323 29882
rect 23013 29824 23018 29880
rect 23074 29824 28262 29880
rect 28318 29824 28323 29880
rect 23013 29822 28323 29824
rect 23013 29819 23079 29822
rect 28257 29819 28323 29822
rect 19568 29408 19888 29409
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 29085 29202 29151 29205
rect 34145 29202 34211 29205
rect 29085 29200 34211 29202
rect 29085 29144 29090 29200
rect 29146 29144 34150 29200
rect 34206 29144 34211 29200
rect 29085 29142 34211 29144
rect 29085 29139 29151 29142
rect 34145 29139 34211 29142
rect 22829 28930 22895 28933
rect 28441 28930 28507 28933
rect 28901 28930 28967 28933
rect 22829 28928 28967 28930
rect 22829 28872 22834 28928
rect 22890 28872 28446 28928
rect 28502 28872 28906 28928
rect 28962 28872 28967 28928
rect 22829 28870 28967 28872
rect 22829 28867 22895 28870
rect 28441 28867 28507 28870
rect 28901 28867 28967 28870
rect 4208 28864 4528 28865
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 30925 28658 30991 28661
rect 33961 28658 34027 28661
rect 30925 28656 34027 28658
rect 30925 28600 30930 28656
rect 30986 28600 33966 28656
rect 34022 28600 34027 28656
rect 30925 28598 34027 28600
rect 30925 28595 30991 28598
rect 33961 28595 34027 28598
rect 28073 28522 28139 28525
rect 32029 28522 32095 28525
rect 28073 28520 32095 28522
rect 28073 28464 28078 28520
rect 28134 28464 32034 28520
rect 32090 28464 32095 28520
rect 28073 28462 32095 28464
rect 28073 28459 28139 28462
rect 32029 28459 32095 28462
rect 31109 28386 31175 28389
rect 32949 28386 33015 28389
rect 33409 28386 33475 28389
rect 31109 28384 33475 28386
rect 31109 28328 31114 28384
rect 31170 28328 32954 28384
rect 33010 28328 33414 28384
rect 33470 28328 33475 28384
rect 31109 28326 33475 28328
rect 31109 28323 31175 28326
rect 32949 28323 33015 28326
rect 33409 28323 33475 28326
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 29177 28248 29243 28253
rect 29177 28192 29182 28248
rect 29238 28192 29243 28248
rect 29177 28187 29243 28192
rect 32121 28250 32187 28253
rect 32673 28250 32739 28253
rect 32121 28248 32739 28250
rect 32121 28192 32126 28248
rect 32182 28192 32678 28248
rect 32734 28192 32739 28248
rect 32121 28190 32739 28192
rect 32121 28187 32187 28190
rect 32673 28187 32739 28190
rect 29180 27981 29240 28187
rect 31845 28114 31911 28117
rect 33225 28114 33291 28117
rect 31845 28112 33291 28114
rect 31845 28056 31850 28112
rect 31906 28056 33230 28112
rect 33286 28056 33291 28112
rect 31845 28054 33291 28056
rect 31845 28051 31911 28054
rect 33225 28051 33291 28054
rect 29177 27976 29243 27981
rect 29177 27920 29182 27976
rect 29238 27920 29243 27976
rect 29177 27915 29243 27920
rect 29361 27978 29427 27981
rect 33685 27978 33751 27981
rect 34789 27978 34855 27981
rect 29361 27976 34855 27978
rect 29361 27920 29366 27976
rect 29422 27920 33690 27976
rect 33746 27920 34794 27976
rect 34850 27920 34855 27976
rect 29361 27918 34855 27920
rect 29361 27915 29427 27918
rect 33685 27915 33751 27918
rect 34789 27915 34855 27918
rect 27429 27842 27495 27845
rect 28441 27842 28507 27845
rect 27429 27840 28507 27842
rect 27429 27784 27434 27840
rect 27490 27784 28446 27840
rect 28502 27784 28507 27840
rect 27429 27782 28507 27784
rect 27429 27779 27495 27782
rect 28441 27779 28507 27782
rect 28993 27842 29059 27845
rect 29637 27842 29703 27845
rect 28993 27840 29703 27842
rect 28993 27784 28998 27840
rect 29054 27784 29642 27840
rect 29698 27784 29703 27840
rect 28993 27782 29703 27784
rect 28993 27779 29059 27782
rect 29637 27779 29703 27782
rect 30833 27842 30899 27845
rect 32581 27842 32647 27845
rect 30833 27840 32647 27842
rect 30833 27784 30838 27840
rect 30894 27784 32586 27840
rect 32642 27784 32647 27840
rect 30833 27782 32647 27784
rect 30833 27779 30899 27782
rect 32581 27779 32647 27782
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 27889 27706 27955 27709
rect 28441 27706 28507 27709
rect 27889 27704 28507 27706
rect 27889 27648 27894 27704
rect 27950 27648 28446 27704
rect 28502 27648 28507 27704
rect 27889 27646 28507 27648
rect 27889 27643 27955 27646
rect 28441 27643 28507 27646
rect 29637 27706 29703 27709
rect 31937 27706 32003 27709
rect 32213 27706 32279 27709
rect 29637 27704 31770 27706
rect 29637 27648 29642 27704
rect 29698 27648 31770 27704
rect 29637 27646 31770 27648
rect 29637 27643 29703 27646
rect 28073 27570 28139 27573
rect 31477 27570 31543 27573
rect 28073 27568 31543 27570
rect 28073 27512 28078 27568
rect 28134 27512 31482 27568
rect 31538 27512 31543 27568
rect 28073 27510 31543 27512
rect 28073 27507 28139 27510
rect 31477 27507 31543 27510
rect 20161 27434 20227 27437
rect 20713 27434 20779 27437
rect 20161 27432 20779 27434
rect 20161 27376 20166 27432
rect 20222 27376 20718 27432
rect 20774 27376 20779 27432
rect 20161 27374 20779 27376
rect 20161 27371 20227 27374
rect 20713 27371 20779 27374
rect 30005 27434 30071 27437
rect 31710 27434 31770 27646
rect 31937 27704 32279 27706
rect 31937 27648 31942 27704
rect 31998 27648 32218 27704
rect 32274 27648 32279 27704
rect 31937 27646 32279 27648
rect 31937 27643 32003 27646
rect 32213 27643 32279 27646
rect 31845 27570 31911 27573
rect 36077 27570 36143 27573
rect 36353 27570 36419 27573
rect 31845 27568 36419 27570
rect 31845 27512 31850 27568
rect 31906 27512 36082 27568
rect 36138 27512 36358 27568
rect 36414 27512 36419 27568
rect 31845 27510 36419 27512
rect 31845 27507 31911 27510
rect 36077 27507 36143 27510
rect 36353 27507 36419 27510
rect 32397 27434 32463 27437
rect 30005 27432 31540 27434
rect 30005 27376 30010 27432
rect 30066 27376 31540 27432
rect 30005 27374 31540 27376
rect 31710 27432 32463 27434
rect 31710 27376 32402 27432
rect 32458 27376 32463 27432
rect 31710 27374 32463 27376
rect 30005 27371 30071 27374
rect 31480 27301 31540 27374
rect 32397 27371 32463 27374
rect 31477 27296 31543 27301
rect 31477 27240 31482 27296
rect 31538 27240 31543 27296
rect 31477 27235 31543 27240
rect 31845 27298 31911 27301
rect 33317 27298 33383 27301
rect 31845 27296 33383 27298
rect 31845 27240 31850 27296
rect 31906 27240 33322 27296
rect 33378 27240 33383 27296
rect 31845 27238 33383 27240
rect 31845 27235 31911 27238
rect 33317 27235 33383 27238
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 27167 19888 27168
rect 20437 27162 20503 27165
rect 25405 27162 25471 27165
rect 20118 27160 25471 27162
rect 20118 27104 20442 27160
rect 20498 27104 25410 27160
rect 25466 27104 25471 27160
rect 20118 27102 25471 27104
rect 18689 27026 18755 27029
rect 20118 27026 20178 27102
rect 20437 27099 20503 27102
rect 25405 27099 25471 27102
rect 25681 27162 25747 27165
rect 35709 27162 35775 27165
rect 25681 27160 35775 27162
rect 25681 27104 25686 27160
rect 25742 27104 35714 27160
rect 35770 27104 35775 27160
rect 25681 27102 35775 27104
rect 25681 27099 25747 27102
rect 35709 27099 35775 27102
rect 22369 27026 22435 27029
rect 25313 27026 25379 27029
rect 27429 27026 27495 27029
rect 18689 27024 20178 27026
rect 18689 26968 18694 27024
rect 18750 26968 20178 27024
rect 18689 26966 20178 26968
rect 20302 27024 27495 27026
rect 20302 26968 22374 27024
rect 22430 26968 25318 27024
rect 25374 26968 27434 27024
rect 27490 26968 27495 27024
rect 20302 26966 27495 26968
rect 18689 26963 18755 26966
rect 19517 26890 19583 26893
rect 20302 26890 20362 26966
rect 22369 26963 22435 26966
rect 25313 26963 25379 26966
rect 27429 26963 27495 26966
rect 31385 27026 31451 27029
rect 32029 27026 32095 27029
rect 36445 27026 36511 27029
rect 31385 27024 36511 27026
rect 31385 26968 31390 27024
rect 31446 26968 32034 27024
rect 32090 26968 36450 27024
rect 36506 26968 36511 27024
rect 31385 26966 36511 26968
rect 31385 26963 31451 26966
rect 32029 26963 32095 26966
rect 36445 26963 36511 26966
rect 19517 26888 20362 26890
rect 19517 26832 19522 26888
rect 19578 26832 20362 26888
rect 19517 26830 20362 26832
rect 28073 26890 28139 26893
rect 32489 26890 32555 26893
rect 28073 26888 32555 26890
rect 28073 26832 28078 26888
rect 28134 26832 32494 26888
rect 32550 26832 32555 26888
rect 28073 26830 32555 26832
rect 19517 26827 19583 26830
rect 28073 26827 28139 26830
rect 32489 26827 32555 26830
rect 20161 26754 20227 26757
rect 28809 26754 28875 26757
rect 20161 26752 28875 26754
rect 20161 26696 20166 26752
rect 20222 26696 28814 26752
rect 28870 26696 28875 26752
rect 20161 26694 28875 26696
rect 20161 26691 20227 26694
rect 28809 26691 28875 26694
rect 29637 26754 29703 26757
rect 33777 26754 33843 26757
rect 29637 26752 33843 26754
rect 29637 26696 29642 26752
rect 29698 26696 33782 26752
rect 33838 26696 33843 26752
rect 29637 26694 33843 26696
rect 29637 26691 29703 26694
rect 33777 26691 33843 26694
rect 4208 26688 4528 26689
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 30097 26618 30163 26621
rect 32857 26618 32923 26621
rect 30097 26616 32923 26618
rect 30097 26560 30102 26616
rect 30158 26560 32862 26616
rect 32918 26560 32923 26616
rect 30097 26558 32923 26560
rect 30097 26555 30163 26558
rect 32857 26555 32923 26558
rect 35341 26618 35407 26621
rect 35893 26618 35959 26621
rect 35341 26616 35959 26618
rect 35341 26560 35346 26616
rect 35402 26560 35898 26616
rect 35954 26560 35959 26616
rect 35341 26558 35959 26560
rect 35341 26555 35407 26558
rect 35893 26555 35959 26558
rect 27061 26482 27127 26485
rect 33593 26482 33659 26485
rect 27061 26480 33659 26482
rect 27061 26424 27066 26480
rect 27122 26424 33598 26480
rect 33654 26424 33659 26480
rect 27061 26422 33659 26424
rect 27061 26419 27127 26422
rect 33593 26419 33659 26422
rect 30005 26346 30071 26349
rect 34053 26346 34119 26349
rect 30005 26344 34119 26346
rect 30005 26288 30010 26344
rect 30066 26288 34058 26344
rect 34114 26288 34119 26344
rect 30005 26286 34119 26288
rect 30005 26283 30071 26286
rect 34053 26283 34119 26286
rect 30925 26212 30991 26213
rect 30925 26210 30972 26212
rect 30880 26208 30972 26210
rect 30880 26152 30930 26208
rect 30880 26150 30972 26152
rect 30925 26148 30972 26150
rect 31036 26148 31042 26212
rect 30925 26147 30991 26148
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 25865 25802 25931 25805
rect 28257 25802 28323 25805
rect 25865 25800 28323 25802
rect 25865 25744 25870 25800
rect 25926 25744 28262 25800
rect 28318 25744 28323 25800
rect 25865 25742 28323 25744
rect 25865 25739 25931 25742
rect 28257 25739 28323 25742
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 30925 25256 30991 25261
rect 30925 25200 30930 25256
rect 30986 25200 30991 25256
rect 30925 25195 30991 25200
rect 19568 25056 19888 25057
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 30741 24986 30807 24989
rect 30928 24986 30988 25195
rect 30741 24984 30988 24986
rect 30741 24928 30746 24984
rect 30802 24928 30988 24984
rect 30741 24926 30988 24928
rect 30741 24923 30807 24926
rect 20529 24850 20595 24853
rect 26233 24850 26299 24853
rect 20529 24848 26299 24850
rect 20529 24792 20534 24848
rect 20590 24792 26238 24848
rect 26294 24792 26299 24848
rect 20529 24790 26299 24792
rect 20529 24787 20595 24790
rect 26233 24787 26299 24790
rect 21817 24578 21883 24581
rect 22185 24578 22251 24581
rect 21817 24576 22251 24578
rect 21817 24520 21822 24576
rect 21878 24520 22190 24576
rect 22246 24520 22251 24576
rect 21817 24518 22251 24520
rect 21817 24515 21883 24518
rect 22185 24515 22251 24518
rect 22737 24578 22803 24581
rect 26417 24578 26483 24581
rect 22737 24576 26483 24578
rect 22737 24520 22742 24576
rect 22798 24520 26422 24576
rect 26478 24520 26483 24576
rect 22737 24518 26483 24520
rect 22737 24515 22803 24518
rect 26417 24515 26483 24518
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 24447 35248 24448
rect 20437 24306 20503 24309
rect 24209 24306 24275 24309
rect 20437 24304 24275 24306
rect 20437 24248 20442 24304
rect 20498 24248 24214 24304
rect 24270 24248 24275 24304
rect 20437 24246 24275 24248
rect 20437 24243 20503 24246
rect 24209 24243 24275 24246
rect 24393 24306 24459 24309
rect 27981 24306 28047 24309
rect 24393 24304 28047 24306
rect 24393 24248 24398 24304
rect 24454 24248 27986 24304
rect 28042 24248 28047 24304
rect 24393 24246 28047 24248
rect 24393 24243 24459 24246
rect 27981 24243 28047 24246
rect 11605 24170 11671 24173
rect 15009 24170 15075 24173
rect 11605 24168 15075 24170
rect 11605 24112 11610 24168
rect 11666 24112 15014 24168
rect 15070 24112 15075 24168
rect 11605 24110 15075 24112
rect 11605 24107 11671 24110
rect 15009 24107 15075 24110
rect 20437 24170 20503 24173
rect 24945 24170 25011 24173
rect 20437 24168 25011 24170
rect 20437 24112 20442 24168
rect 20498 24112 24950 24168
rect 25006 24112 25011 24168
rect 20437 24110 25011 24112
rect 20437 24107 20503 24110
rect 24945 24107 25011 24110
rect 21173 24034 21239 24037
rect 24301 24034 24367 24037
rect 21173 24032 24367 24034
rect 21173 23976 21178 24032
rect 21234 23976 24306 24032
rect 24362 23976 24367 24032
rect 21173 23974 24367 23976
rect 21173 23971 21239 23974
rect 24301 23971 24367 23974
rect 19568 23968 19888 23969
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 22093 23898 22159 23901
rect 22737 23898 22803 23901
rect 28165 23898 28231 23901
rect 22093 23896 28231 23898
rect 22093 23840 22098 23896
rect 22154 23840 22742 23896
rect 22798 23840 28170 23896
rect 28226 23840 28231 23896
rect 22093 23838 28231 23840
rect 22093 23835 22159 23838
rect 22737 23835 22803 23838
rect 28165 23835 28231 23838
rect 21081 23626 21147 23629
rect 22461 23626 22527 23629
rect 21081 23624 22527 23626
rect 21081 23568 21086 23624
rect 21142 23568 22466 23624
rect 22522 23568 22527 23624
rect 21081 23566 22527 23568
rect 21081 23563 21147 23566
rect 22461 23563 22527 23566
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 21541 23354 21607 23357
rect 29361 23354 29427 23357
rect 21541 23352 29427 23354
rect 21541 23296 21546 23352
rect 21602 23296 29366 23352
rect 29422 23296 29427 23352
rect 21541 23294 29427 23296
rect 21541 23291 21607 23294
rect 29361 23291 29427 23294
rect 34513 23218 34579 23221
rect 39200 23218 40000 23248
rect 34513 23216 40000 23218
rect 34513 23160 34518 23216
rect 34574 23160 40000 23216
rect 34513 23158 40000 23160
rect 34513 23155 34579 23158
rect 39200 23128 40000 23158
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 15837 21994 15903 21997
rect 20437 21994 20503 21997
rect 15837 21992 20503 21994
rect 15837 21936 15842 21992
rect 15898 21936 20442 21992
rect 20498 21936 20503 21992
rect 15837 21934 20503 21936
rect 15837 21931 15903 21934
rect 20437 21931 20503 21934
rect 0 21858 800 21888
rect 1393 21858 1459 21861
rect 0 21856 1459 21858
rect 0 21800 1398 21856
rect 1454 21800 1459 21856
rect 0 21798 1459 21800
rect 0 21768 800 21798
rect 1393 21795 1459 21798
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 21727 19888 21728
rect 25865 21722 25931 21725
rect 30741 21722 30807 21725
rect 25865 21720 30807 21722
rect 25865 21664 25870 21720
rect 25926 21664 30746 21720
rect 30802 21664 30807 21720
rect 25865 21662 30807 21664
rect 25865 21659 25931 21662
rect 30741 21659 30807 21662
rect 15377 21586 15443 21589
rect 18321 21586 18387 21589
rect 18597 21586 18663 21589
rect 15377 21584 18663 21586
rect 15377 21528 15382 21584
rect 15438 21528 18326 21584
rect 18382 21528 18602 21584
rect 18658 21528 18663 21584
rect 15377 21526 18663 21528
rect 15377 21523 15443 21526
rect 18321 21523 18387 21526
rect 18597 21523 18663 21526
rect 22001 21586 22067 21589
rect 24301 21586 24367 21589
rect 22001 21584 24367 21586
rect 22001 21528 22006 21584
rect 22062 21528 24306 21584
rect 24362 21528 24367 21584
rect 22001 21526 24367 21528
rect 22001 21523 22067 21526
rect 24301 21523 24367 21526
rect 30557 21586 30623 21589
rect 38101 21586 38167 21589
rect 30557 21584 38167 21586
rect 30557 21528 30562 21584
rect 30618 21528 38106 21584
rect 38162 21528 38167 21584
rect 30557 21526 38167 21528
rect 30557 21523 30623 21526
rect 38101 21523 38167 21526
rect 4208 21248 4528 21249
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 27429 20634 27495 20637
rect 27981 20634 28047 20637
rect 27429 20632 28047 20634
rect 27429 20576 27434 20632
rect 27490 20576 27986 20632
rect 28042 20576 28047 20632
rect 27429 20574 28047 20576
rect 27429 20571 27495 20574
rect 27981 20571 28047 20574
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 23657 20090 23723 20093
rect 26049 20090 26115 20093
rect 23657 20088 26115 20090
rect 23657 20032 23662 20088
rect 23718 20032 26054 20088
rect 26110 20032 26115 20088
rect 23657 20030 26115 20032
rect 23657 20027 23723 20030
rect 26049 20027 26115 20030
rect 23473 19818 23539 19821
rect 27981 19818 28047 19821
rect 23473 19816 28047 19818
rect 23473 19760 23478 19816
rect 23534 19760 27986 19816
rect 28042 19760 28047 19816
rect 23473 19758 28047 19760
rect 23473 19755 23539 19758
rect 27981 19755 28047 19758
rect 27337 19682 27403 19685
rect 28901 19682 28967 19685
rect 27337 19680 28967 19682
rect 27337 19624 27342 19680
rect 27398 19624 28906 19680
rect 28962 19624 28967 19680
rect 27337 19622 28967 19624
rect 27337 19619 27403 19622
rect 28901 19619 28967 19622
rect 19568 19616 19888 19617
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 10409 19546 10475 19549
rect 12341 19546 12407 19549
rect 10409 19544 12407 19546
rect 10409 19488 10414 19544
rect 10470 19488 12346 19544
rect 12402 19488 12407 19544
rect 10409 19486 12407 19488
rect 10409 19483 10475 19486
rect 12341 19483 12407 19486
rect 20161 19546 20227 19549
rect 20345 19546 20411 19549
rect 20161 19544 20411 19546
rect 20161 19488 20166 19544
rect 20222 19488 20350 19544
rect 20406 19488 20411 19544
rect 20161 19486 20411 19488
rect 20161 19483 20227 19486
rect 20345 19483 20411 19486
rect 9673 19410 9739 19413
rect 10593 19410 10659 19413
rect 9673 19408 10659 19410
rect 9673 19352 9678 19408
rect 9734 19352 10598 19408
rect 10654 19352 10659 19408
rect 9673 19350 10659 19352
rect 9673 19347 9739 19350
rect 10593 19347 10659 19350
rect 19793 19410 19859 19413
rect 23657 19410 23723 19413
rect 19793 19408 23723 19410
rect 19793 19352 19798 19408
rect 19854 19352 23662 19408
rect 23718 19352 23723 19408
rect 19793 19350 23723 19352
rect 19793 19347 19859 19350
rect 23657 19347 23723 19350
rect 29637 19410 29703 19413
rect 30373 19410 30439 19413
rect 29637 19408 30439 19410
rect 29637 19352 29642 19408
rect 29698 19352 30378 19408
rect 30434 19352 30439 19408
rect 29637 19350 30439 19352
rect 29637 19347 29703 19350
rect 30373 19347 30439 19350
rect 19793 19274 19859 19277
rect 20529 19274 20595 19277
rect 19793 19272 20595 19274
rect 19793 19216 19798 19272
rect 19854 19216 20534 19272
rect 20590 19216 20595 19272
rect 19793 19214 20595 19216
rect 19793 19211 19859 19214
rect 20529 19211 20595 19214
rect 25773 19274 25839 19277
rect 28717 19274 28783 19277
rect 25773 19272 28783 19274
rect 25773 19216 25778 19272
rect 25834 19216 28722 19272
rect 28778 19216 28783 19272
rect 25773 19214 28783 19216
rect 25773 19211 25839 19214
rect 28717 19211 28783 19214
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 19007 35248 19008
rect 19701 18866 19767 18869
rect 24301 18866 24367 18869
rect 19701 18864 24367 18866
rect 19701 18808 19706 18864
rect 19762 18808 24306 18864
rect 24362 18808 24367 18864
rect 19701 18806 24367 18808
rect 19701 18803 19767 18806
rect 24301 18803 24367 18806
rect 15285 18730 15351 18733
rect 18413 18730 18479 18733
rect 15285 18728 18479 18730
rect 15285 18672 15290 18728
rect 15346 18672 18418 18728
rect 18474 18672 18479 18728
rect 15285 18670 18479 18672
rect 15285 18667 15351 18670
rect 18413 18667 18479 18670
rect 19568 18528 19888 18529
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 16287 19888 16288
rect 4208 15808 4528 15809
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 21817 14378 21883 14381
rect 22737 14378 22803 14381
rect 21817 14376 22803 14378
rect 21817 14320 21822 14376
rect 21878 14320 22742 14376
rect 22798 14320 22803 14376
rect 21817 14318 22803 14320
rect 21817 14315 21883 14318
rect 22737 14315 22803 14318
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 13567 35248 13568
rect 14733 13290 14799 13293
rect 15745 13290 15811 13293
rect 14733 13288 15811 13290
rect 14733 13232 14738 13288
rect 14794 13232 15750 13288
rect 15806 13232 15811 13288
rect 14733 13230 15811 13232
rect 14733 13227 14799 13230
rect 15745 13227 15811 13230
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 9949 12474 10015 12477
rect 17217 12474 17283 12477
rect 9949 12472 17283 12474
rect 9949 12416 9954 12472
rect 10010 12416 17222 12472
rect 17278 12416 17283 12472
rect 9949 12414 17283 12416
rect 9949 12411 10015 12414
rect 17217 12411 17283 12414
rect 38009 12338 38075 12341
rect 39200 12338 40000 12368
rect 38009 12336 40000 12338
rect 38009 12280 38014 12336
rect 38070 12280 40000 12336
rect 38009 12278 40000 12280
rect 38009 12275 38075 12278
rect 39200 12248 40000 12278
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 0 10978 800 11008
rect 1577 10978 1643 10981
rect 0 10976 1643 10978
rect 0 10920 1582 10976
rect 1638 10920 1643 10976
rect 0 10918 1643 10920
rect 0 10888 800 10918
rect 1577 10915 1643 10918
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 4208 10368 4528 10369
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 8127 35248 8128
rect 19568 7648 19888 7649
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 5407 19888 5408
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2687 35248 2688
rect 19568 2208 19888 2209
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
rect 38009 1458 38075 1461
rect 39200 1458 40000 1488
rect 38009 1456 40000 1458
rect 38009 1400 38014 1456
rect 38070 1400 40000 1456
rect 38009 1398 40000 1400
rect 38009 1395 38075 1398
rect 39200 1368 40000 1398
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 30788 31920 30852 31924
rect 30788 31864 30802 31920
rect 30802 31864 30852 31920
rect 30788 31860 30852 31864
rect 30972 31588 31036 31652
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 30788 31512 30852 31516
rect 30788 31456 30802 31512
rect 30802 31456 30852 31512
rect 30788 31452 30852 31456
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 30972 26208 31036 26212
rect 30972 26152 30986 26208
rect 30986 26152 31036 26208
rect 30972 26148 31036 26152
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36212 4528 36416
rect 4208 35976 4250 36212
rect 4486 35976 4528 36212
rect 4208 35392 4528 35976
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5576 4528 5952
rect 4208 5340 4250 5576
rect 4486 5340 4528 5576
rect 4208 4928 4528 5340
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36212 35248 36416
rect 34928 35976 34970 36212
rect 35206 35976 35248 36212
rect 34928 35392 35248 35976
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 30787 31924 30853 31925
rect 30787 31860 30788 31924
rect 30852 31860 30853 31924
rect 30787 31859 30853 31860
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 30790 31517 30850 31859
rect 30971 31652 31037 31653
rect 30971 31588 30972 31652
rect 31036 31588 31037 31652
rect 30971 31587 31037 31588
rect 30787 31516 30853 31517
rect 30787 31452 30788 31516
rect 30852 31452 30853 31516
rect 30787 31451 30853 31452
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 30974 26213 31034 31587
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 30971 26212 31037 26213
rect 30971 26148 30972 26212
rect 31036 26148 31037 26212
rect 30971 26147 31037 26148
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20894 19888 21728
rect 19568 20704 19610 20894
rect 19846 20704 19888 20894
rect 19568 20640 19576 20704
rect 19640 20640 19656 20658
rect 19720 20640 19736 20658
rect 19800 20640 19816 20658
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5576 35248 5952
rect 34928 5340 34970 5576
rect 35206 5340 35248 5576
rect 34928 4928 35248 5340
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
<< via4 >>
rect 4250 35976 4486 36212
rect 4250 5340 4486 5576
rect 34970 35976 35206 36212
rect 19610 20704 19846 20894
rect 19610 20658 19640 20704
rect 19640 20658 19656 20704
rect 19656 20658 19720 20704
rect 19720 20658 19736 20704
rect 19736 20658 19800 20704
rect 19800 20658 19816 20704
rect 19816 20658 19846 20704
rect 34970 5340 35206 5576
<< metal5 >>
rect 1104 36212 38824 36254
rect 1104 35976 4250 36212
rect 4486 35976 34970 36212
rect 35206 35976 38824 36212
rect 1104 35934 38824 35976
rect 1104 20894 38824 20936
rect 1104 20658 19610 20894
rect 19846 20658 38824 20894
rect 1104 20616 38824 20658
rect 1104 5576 38824 5618
rect 1104 5340 4250 5576
rect 4486 5340 34970 5576
rect 35206 5340 38824 5576
rect 1104 5298 38824 5340
use sky130_fd_sc_hd__diode_2  ANTENNA_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 17388 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1656 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2760 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_29
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_41
timestamp 1644511149
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_57
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_69
timestamp 1644511149
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1644511149
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_85
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_97 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_104
timestamp 1644511149
transform 1 0 10672 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_113
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1644511149
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1644511149
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_153
timestamp 1644511149
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1644511149
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_169
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_181
timestamp 1644511149
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1644511149
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_197
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_209
timestamp 1644511149
transform 1 0 20332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_217 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21068 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_225
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_237
timestamp 1644511149
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1644511149
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_253
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_265
timestamp 1644511149
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1644511149
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_281
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_293
timestamp 1644511149
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1644511149
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_309
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_321
timestamp 1644511149
transform 1 0 30636 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_332
timestamp 1644511149
transform 1 0 31648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_337
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_349
timestamp 1644511149
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1644511149
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_365
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_377
timestamp 1644511149
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 1644511149
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_393
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_403
timestamp 1644511149
transform 1 0 38180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1644511149
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1644511149
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1644511149
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1644511149
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1644511149
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_69
timestamp 1644511149
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_81
timestamp 1644511149
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_93
timestamp 1644511149
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1644511149
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1644511149
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_113
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_125
timestamp 1644511149
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_137
timestamp 1644511149
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_149
timestamp 1644511149
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1644511149
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1644511149
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_169
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_181
timestamp 1644511149
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_193
timestamp 1644511149
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_205
timestamp 1644511149
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1644511149
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1644511149
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_225
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_237
timestamp 1644511149
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_249
timestamp 1644511149
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_261
timestamp 1644511149
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1644511149
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1644511149
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_281
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_293
timestamp 1644511149
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_305
timestamp 1644511149
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_317
timestamp 1644511149
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1644511149
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1644511149
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_337
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_349
timestamp 1644511149
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_361
timestamp 1644511149
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_373
timestamp 1644511149
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1644511149
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1644511149
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_393
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp 1644511149
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1644511149
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1644511149
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_29
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_41
timestamp 1644511149
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_53
timestamp 1644511149
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_65
timestamp 1644511149
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1644511149
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1644511149
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_97
timestamp 1644511149
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_109
timestamp 1644511149
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_121
timestamp 1644511149
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1644511149
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1644511149
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_153
timestamp 1644511149
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_165
timestamp 1644511149
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_177
timestamp 1644511149
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1644511149
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1644511149
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_197
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_209
timestamp 1644511149
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_221
timestamp 1644511149
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_233
timestamp 1644511149
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1644511149
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1644511149
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_265
timestamp 1644511149
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_277
timestamp 1644511149
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_289
timestamp 1644511149
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1644511149
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1644511149
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_309
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_321
timestamp 1644511149
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_333
timestamp 1644511149
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_345
timestamp 1644511149
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1644511149
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1644511149
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_377
timestamp 1644511149
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_389
timestamp 1644511149
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_401
timestamp 1644511149
transform 1 0 37996 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1644511149
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1644511149
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1644511149
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1644511149
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1644511149
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_57
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_69
timestamp 1644511149
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_81
timestamp 1644511149
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_93
timestamp 1644511149
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1644511149
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1644511149
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_125
timestamp 1644511149
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_137
timestamp 1644511149
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_149
timestamp 1644511149
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1644511149
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1644511149
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_181
timestamp 1644511149
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_193
timestamp 1644511149
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_205
timestamp 1644511149
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1644511149
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1644511149
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_225
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_237
timestamp 1644511149
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_249
timestamp 1644511149
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_261
timestamp 1644511149
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1644511149
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1644511149
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_293
timestamp 1644511149
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_305
timestamp 1644511149
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_317
timestamp 1644511149
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1644511149
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1644511149
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_337
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_349
timestamp 1644511149
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_361
timestamp 1644511149
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_373
timestamp 1644511149
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1644511149
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1644511149
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_393
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 1644511149
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1644511149
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1644511149
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_29
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_41
timestamp 1644511149
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_53
timestamp 1644511149
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_65
timestamp 1644511149
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1644511149
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1644511149
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_97
timestamp 1644511149
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_109
timestamp 1644511149
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_121
timestamp 1644511149
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1644511149
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1644511149
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_165
timestamp 1644511149
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_177
timestamp 1644511149
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1644511149
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1644511149
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_209
timestamp 1644511149
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_221
timestamp 1644511149
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_233
timestamp 1644511149
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1644511149
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1644511149
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_265
timestamp 1644511149
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_277
timestamp 1644511149
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_289
timestamp 1644511149
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1644511149
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1644511149
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_309
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_321
timestamp 1644511149
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_333
timestamp 1644511149
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_345
timestamp 1644511149
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1644511149
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1644511149
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_365
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_377
timestamp 1644511149
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_389
timestamp 1644511149
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_401
timestamp 1644511149
transform 1 0 37996 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1644511149
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1644511149
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1644511149
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1644511149
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1644511149
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1644511149
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1644511149
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1644511149
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1644511149
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_181
timestamp 1644511149
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_193
timestamp 1644511149
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_205
timestamp 1644511149
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1644511149
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1644511149
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_237
timestamp 1644511149
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_249
timestamp 1644511149
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_261
timestamp 1644511149
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1644511149
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1644511149
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_305
timestamp 1644511149
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_317
timestamp 1644511149
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1644511149
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1644511149
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_349
timestamp 1644511149
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_361
timestamp 1644511149
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_373
timestamp 1644511149
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1644511149
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1644511149
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_393
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_405
timestamp 1644511149
transform 1 0 38364 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1644511149
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1644511149
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1644511149
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1644511149
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1644511149
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_177
timestamp 1644511149
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1644511149
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_209
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_221
timestamp 1644511149
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_233
timestamp 1644511149
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1644511149
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1644511149
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1644511149
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_277
timestamp 1644511149
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_289
timestamp 1644511149
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1644511149
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_321
timestamp 1644511149
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_333
timestamp 1644511149
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_345
timestamp 1644511149
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1644511149
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_365
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_377
timestamp 1644511149
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_389
timestamp 1644511149
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_401
timestamp 1644511149
transform 1 0 37996 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1644511149
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1644511149
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1644511149
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1644511149
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1644511149
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1644511149
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_193
timestamp 1644511149
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_205
timestamp 1644511149
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1644511149
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_249
timestamp 1644511149
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_261
timestamp 1644511149
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1644511149
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1644511149
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_317
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1644511149
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1644511149
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_361
timestamp 1644511149
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_373
timestamp 1644511149
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1644511149
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1644511149
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_405
timestamp 1644511149
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1644511149
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1644511149
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1644511149
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_91
timestamp 1644511149
transform 1 0 9476 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_103
timestamp 1644511149
transform 1 0 10580 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_115
timestamp 1644511149
transform 1 0 11684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_127
timestamp 1644511149
transform 1 0 12788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_165
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_177
timestamp 1644511149
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1644511149
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_209
timestamp 1644511149
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_221
timestamp 1644511149
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_233
timestamp 1644511149
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1644511149
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1644511149
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_265
timestamp 1644511149
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_277
timestamp 1644511149
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_289
timestamp 1644511149
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1644511149
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_321
timestamp 1644511149
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_333
timestamp 1644511149
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_345
timestamp 1644511149
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1644511149
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1644511149
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_377
timestamp 1644511149
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_389
timestamp 1644511149
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_401
timestamp 1644511149
transform 1 0 37996 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1644511149
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1644511149
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1644511149
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1644511149
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_97
timestamp 1644511149
transform 1 0 10028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_109
timestamp 1644511149
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_180
timestamp 1644511149
transform 1 0 17664 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_192
timestamp 1644511149
transform 1 0 18768 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_204
timestamp 1644511149
transform 1 0 19872 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_216
timestamp 1644511149
transform 1 0 20976 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_237
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_261
timestamp 1644511149
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1644511149
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_293
timestamp 1644511149
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_305
timestamp 1644511149
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_317
timestamp 1644511149
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1644511149
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1644511149
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_349
timestamp 1644511149
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_361
timestamp 1644511149
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_373
timestamp 1644511149
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1644511149
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1644511149
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1644511149
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1644511149
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1644511149
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_107
timestamp 1644511149
transform 1 0 10948 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_116
timestamp 1644511149
transform 1 0 11776 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_123
timestamp 1644511149
transform 1 0 12420 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_135
timestamp 1644511149
transform 1 0 13524 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_165
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_173
timestamp 1644511149
transform 1 0 17020 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_191
timestamp 1644511149
transform 1 0 18676 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_209
timestamp 1644511149
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_221
timestamp 1644511149
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_233
timestamp 1644511149
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1644511149
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1644511149
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_265
timestamp 1644511149
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_277
timestamp 1644511149
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_289
timestamp 1644511149
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1644511149
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1644511149
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_321
timestamp 1644511149
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_333
timestamp 1644511149
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_345
timestamp 1644511149
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1644511149
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1644511149
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_365
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_377
timestamp 1644511149
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_389
timestamp 1644511149
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_401
timestamp 1644511149
transform 1 0 37996 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1644511149
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1644511149
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1644511149
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1644511149
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_93
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_100
timestamp 1644511149
transform 1 0 10304 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_107
timestamp 1644511149
transform 1 0 10948 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1644511149
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_131
timestamp 1644511149
transform 1 0 13156 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_143
timestamp 1644511149
transform 1 0 14260 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_147
timestamp 1644511149
transform 1 0 14628 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_164
timestamp 1644511149
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_173
timestamp 1644511149
transform 1 0 17020 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_177
timestamp 1644511149
transform 1 0 17388 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_189
timestamp 1644511149
transform 1 0 18492 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_201
timestamp 1644511149
transform 1 0 19596 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_213
timestamp 1644511149
transform 1 0 20700 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_221
timestamp 1644511149
transform 1 0 21436 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_237
timestamp 1644511149
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_249
timestamp 1644511149
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_261
timestamp 1644511149
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1644511149
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1644511149
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_293
timestamp 1644511149
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_305
timestamp 1644511149
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_317
timestamp 1644511149
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1644511149
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1644511149
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_361
timestamp 1644511149
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_373
timestamp 1644511149
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1644511149
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1644511149
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_405
timestamp 1644511149
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1644511149
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1644511149
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_73
timestamp 1644511149
transform 1 0 7820 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_80
timestamp 1644511149
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_96
timestamp 1644511149
transform 1 0 9936 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_116
timestamp 1644511149
transform 1 0 11776 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_125
timestamp 1644511149
transform 1 0 12604 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_136
timestamp 1644511149
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_157
timestamp 1644511149
transform 1 0 15548 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_166
timestamp 1644511149
transform 1 0 16376 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_173
timestamp 1644511149
transform 1 0 17020 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_181
timestamp 1644511149
transform 1 0 17756 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_191
timestamp 1644511149
transform 1 0 18676 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1644511149
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_202
timestamp 1644511149
transform 1 0 19688 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_206
timestamp 1644511149
transform 1 0 20056 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_212
timestamp 1644511149
transform 1 0 20608 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_219
timestamp 1644511149
transform 1 0 21252 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_227
timestamp 1644511149
transform 1 0 21988 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_231
timestamp 1644511149
transform 1 0 22356 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_238
timestamp 1644511149
transform 1 0 23000 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_250
timestamp 1644511149
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_265
timestamp 1644511149
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_277
timestamp 1644511149
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_289
timestamp 1644511149
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1644511149
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1644511149
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_321
timestamp 1644511149
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_333
timestamp 1644511149
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_345
timestamp 1644511149
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1644511149
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1644511149
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_377
timestamp 1644511149
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_389
timestamp 1644511149
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_401
timestamp 1644511149
transform 1 0 37996 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1644511149
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1644511149
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1644511149
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_65
timestamp 1644511149
transform 1 0 7084 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_82
timestamp 1644511149
transform 1 0 8648 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_89
timestamp 1644511149
transform 1 0 9292 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_101
timestamp 1644511149
transform 1 0 10396 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_108
timestamp 1644511149
transform 1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_119
timestamp 1644511149
transform 1 0 12052 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_131
timestamp 1644511149
transform 1 0 13156 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_149
timestamp 1644511149
transform 1 0 14812 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_156
timestamp 1644511149
transform 1 0 15456 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_160
timestamp 1644511149
transform 1 0 15824 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_164
timestamp 1644511149
transform 1 0 16192 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_174
timestamp 1644511149
transform 1 0 17112 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_13_196
timestamp 1644511149
transform 1 0 19136 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_220
timestamp 1644511149
transform 1 0 21344 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_245
timestamp 1644511149
transform 1 0 23644 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_257
timestamp 1644511149
transform 1 0 24748 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_269
timestamp 1644511149
transform 1 0 25852 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_277
timestamp 1644511149
transform 1 0 26588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_293
timestamp 1644511149
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_305
timestamp 1644511149
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_317
timestamp 1644511149
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1644511149
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1644511149
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_349
timestamp 1644511149
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_361
timestamp 1644511149
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_373
timestamp 1644511149
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1644511149
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1644511149
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1644511149
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1644511149
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_73
timestamp 1644511149
transform 1 0 7820 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_80
timestamp 1644511149
transform 1 0 8464 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_94
timestamp 1644511149
transform 1 0 9752 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_103
timestamp 1644511149
transform 1 0 10580 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_123
timestamp 1644511149
transform 1 0 12420 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_132
timestamp 1644511149
transform 1 0 13248 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_146
timestamp 1644511149
transform 1 0 14536 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_153
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_157
timestamp 1644511149
transform 1 0 15548 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_174
timestamp 1644511149
transform 1 0 17112 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_184
timestamp 1644511149
transform 1 0 18032 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_191
timestamp 1644511149
transform 1 0 18676 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1644511149
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_213
timestamp 1644511149
transform 1 0 20700 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_221
timestamp 1644511149
transform 1 0 21436 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_239
timestamp 1644511149
transform 1 0 23092 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1644511149
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_257
timestamp 1644511149
transform 1 0 24748 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_266
timestamp 1644511149
transform 1 0 25576 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_278
timestamp 1644511149
transform 1 0 26680 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_290
timestamp 1644511149
transform 1 0 27784 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_302
timestamp 1644511149
transform 1 0 28888 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_321
timestamp 1644511149
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_333
timestamp 1644511149
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_345
timestamp 1644511149
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1644511149
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1644511149
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_389
timestamp 1644511149
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_401
timestamp 1644511149
transform 1 0 37996 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1644511149
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1644511149
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1644511149
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1644511149
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_73
timestamp 1644511149
transform 1 0 7820 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_82
timestamp 1644511149
transform 1 0 8648 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_15_94
timestamp 1644511149
transform 1 0 9752 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_100
timestamp 1644511149
transform 1 0 10304 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_108
timestamp 1644511149
transform 1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_121
timestamp 1644511149
transform 1 0 12236 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_129
timestamp 1644511149
transform 1 0 12972 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_146
timestamp 1644511149
transform 1 0 14536 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_156
timestamp 1644511149
transform 1 0 15456 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_163
timestamp 1644511149
transform 1 0 16100 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1644511149
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_177
timestamp 1644511149
transform 1 0 17388 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_189
timestamp 1644511149
transform 1 0 18492 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_197
timestamp 1644511149
transform 1 0 19228 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_204
timestamp 1644511149
transform 1 0 19872 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_214
timestamp 1644511149
transform 1 0 20792 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1644511149
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_230
timestamp 1644511149
transform 1 0 22264 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_239
timestamp 1644511149
transform 1 0 23092 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_251
timestamp 1644511149
transform 1 0 24196 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_258
timestamp 1644511149
transform 1 0 24840 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_266
timestamp 1644511149
transform 1 0 25576 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_276
timestamp 1644511149
transform 1 0 26496 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_293
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_305
timestamp 1644511149
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_317
timestamp 1644511149
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1644511149
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1644511149
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_373
timestamp 1644511149
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1644511149
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1644511149
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_7
timestamp 1644511149
transform 1 0 1748 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_19
timestamp 1644511149
transform 1 0 2852 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1644511149
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_61
timestamp 1644511149
transform 1 0 6716 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_80
timestamp 1644511149
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_101
timestamp 1644511149
transform 1 0 10396 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_121
timestamp 1644511149
transform 1 0 12236 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_129
timestamp 1644511149
transform 1 0 12972 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_136
timestamp 1644511149
transform 1 0 13616 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_149
timestamp 1644511149
transform 1 0 14812 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_157
timestamp 1644511149
transform 1 0 15548 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_166
timestamp 1644511149
transform 1 0 16376 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_186
timestamp 1644511149
transform 1 0 18216 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1644511149
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_200
timestamp 1644511149
transform 1 0 19504 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_212
timestamp 1644511149
transform 1 0 20608 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_229
timestamp 1644511149
transform 1 0 22172 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_241
timestamp 1644511149
transform 1 0 23276 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_248
timestamp 1644511149
transform 1 0 23920 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_261
timestamp 1644511149
transform 1 0 25116 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_286
timestamp 1644511149
transform 1 0 27416 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_298
timestamp 1644511149
transform 1 0 28520 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_306
timestamp 1644511149
transform 1 0 29256 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_321
timestamp 1644511149
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_333
timestamp 1644511149
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_345
timestamp 1644511149
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1644511149
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1644511149
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_377
timestamp 1644511149
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_389
timestamp 1644511149
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_401
timestamp 1644511149
transform 1 0 37996 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1644511149
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1644511149
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1644511149
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1644511149
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1644511149
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_77
timestamp 1644511149
transform 1 0 8188 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_83
timestamp 1644511149
transform 1 0 8740 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_94
timestamp 1644511149
transform 1 0 9752 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_108
timestamp 1644511149
transform 1 0 11040 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_117
timestamp 1644511149
transform 1 0 11868 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_125
timestamp 1644511149
transform 1 0 12604 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_137
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_144
timestamp 1644511149
transform 1 0 14352 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_164
timestamp 1644511149
transform 1 0 16192 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_179
timestamp 1644511149
transform 1 0 17572 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_187
timestamp 1644511149
transform 1 0 18308 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_195
timestamp 1644511149
transform 1 0 19044 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_201
timestamp 1644511149
transform 1 0 19596 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_210
timestamp 1644511149
transform 1 0 20424 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1644511149
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1644511149
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_233
timestamp 1644511149
transform 1 0 22540 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_241
timestamp 1644511149
transform 1 0 23276 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_255
timestamp 1644511149
transform 1 0 24564 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_265
timestamp 1644511149
transform 1 0 25484 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_274
timestamp 1644511149
transform 1 0 26312 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_284
timestamp 1644511149
transform 1 0 27232 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_291
timestamp 1644511149
transform 1 0 27876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_303
timestamp 1644511149
transform 1 0 28980 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_315
timestamp 1644511149
transform 1 0 30084 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_327
timestamp 1644511149
transform 1 0 31188 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1644511149
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_349
timestamp 1644511149
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_361
timestamp 1644511149
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_373
timestamp 1644511149
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1644511149
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1644511149
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1644511149
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1644511149
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1644511149
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_88
timestamp 1644511149
transform 1 0 9200 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_108
timestamp 1644511149
transform 1 0 11040 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_117
timestamp 1644511149
transform 1 0 11868 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_126
timestamp 1644511149
transform 1 0 12696 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1644511149
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_146
timestamp 1644511149
transform 1 0 14536 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_155
timestamp 1644511149
transform 1 0 15364 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_169
timestamp 1644511149
transform 1 0 16652 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_177
timestamp 1644511149
transform 1 0 17388 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_192
timestamp 1644511149
transform 1 0 18768 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_213
timestamp 1644511149
transform 1 0 20700 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_220
timestamp 1644511149
transform 1 0 21344 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_233
timestamp 1644511149
transform 1 0 22540 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_246
timestamp 1644511149
transform 1 0 23736 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_18_263
timestamp 1644511149
transform 1 0 25300 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_278
timestamp 1644511149
transform 1 0 26680 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_287
timestamp 1644511149
transform 1 0 27508 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_299
timestamp 1644511149
transform 1 0 28612 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1644511149
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_321
timestamp 1644511149
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_333
timestamp 1644511149
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_345
timestamp 1644511149
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1644511149
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1644511149
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_377
timestamp 1644511149
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_389
timestamp 1644511149
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_401
timestamp 1644511149
transform 1 0 37996 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1644511149
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1644511149
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1644511149
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1644511149
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_91
timestamp 1644511149
transform 1 0 9476 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_100
timestamp 1644511149
transform 1 0 10304 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_104
timestamp 1644511149
transform 1 0 10672 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_108
timestamp 1644511149
transform 1 0 11040 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_129
timestamp 1644511149
transform 1 0 12972 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_149
timestamp 1644511149
transform 1 0 14812 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_159
timestamp 1644511149
transform 1 0 15732 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1644511149
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_172
timestamp 1644511149
transform 1 0 16928 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_192
timestamp 1644511149
transform 1 0 18768 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_200
timestamp 1644511149
transform 1 0 19504 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_210
timestamp 1644511149
transform 1 0 20424 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1644511149
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_234
timestamp 1644511149
transform 1 0 22632 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_251
timestamp 1644511149
transform 1 0 24196 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_255
timestamp 1644511149
transform 1 0 24564 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_263
timestamp 1644511149
transform 1 0 25300 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_267
timestamp 1644511149
transform 1 0 25668 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_276
timestamp 1644511149
transform 1 0 26496 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_290
timestamp 1644511149
transform 1 0 27784 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_299
timestamp 1644511149
transform 1 0 28612 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_311
timestamp 1644511149
transform 1 0 29716 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_323
timestamp 1644511149
transform 1 0 30820 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1644511149
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_337
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_349
timestamp 1644511149
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_361
timestamp 1644511149
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_373
timestamp 1644511149
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1644511149
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1644511149
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_403
timestamp 1644511149
transform 1 0 38180 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1644511149
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1644511149
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_61
timestamp 1644511149
transform 1 0 6716 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_80
timestamp 1644511149
transform 1 0 8464 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_88
timestamp 1644511149
transform 1 0 9200 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_92
timestamp 1644511149
transform 1 0 9568 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_99
timestamp 1644511149
transform 1 0 10212 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_111
timestamp 1644511149
transform 1 0 11316 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_117
timestamp 1644511149
transform 1 0 11868 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_123
timestamp 1644511149
transform 1 0 12420 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_127
timestamp 1644511149
transform 1 0 12788 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_136
timestamp 1644511149
transform 1 0 13616 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_152
timestamp 1644511149
transform 1 0 15088 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_172
timestamp 1644511149
transform 1 0 16928 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_180
timestamp 1644511149
transform 1 0 17664 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_187
timestamp 1644511149
transform 1 0 18308 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1644511149
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_202
timestamp 1644511149
transform 1 0 19688 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_217
timestamp 1644511149
transform 1 0 21068 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_237
timestamp 1644511149
transform 1 0 22908 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_243
timestamp 1644511149
transform 1 0 23460 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_248
timestamp 1644511149
transform 1 0 23920 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_262
timestamp 1644511149
transform 1 0 25208 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_280
timestamp 1644511149
transform 1 0 26864 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_294
timestamp 1644511149
transform 1 0 28152 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_306
timestamp 1644511149
transform 1 0 29256 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_321
timestamp 1644511149
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_333
timestamp 1644511149
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_345
timestamp 1644511149
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1644511149
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1644511149
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_377
timestamp 1644511149
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_389
timestamp 1644511149
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_401
timestamp 1644511149
transform 1 0 37996 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1644511149
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1644511149
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1644511149
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1644511149
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_77
timestamp 1644511149
transform 1 0 8188 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_86
timestamp 1644511149
transform 1 0 9016 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_97
timestamp 1644511149
transform 1 0 10028 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_104
timestamp 1644511149
transform 1 0 10672 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_116
timestamp 1644511149
transform 1 0 11776 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_124
timestamp 1644511149
transform 1 0 12512 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_137
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_157
timestamp 1644511149
transform 1 0 15548 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_164
timestamp 1644511149
transform 1 0 16192 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_183
timestamp 1644511149
transform 1 0 17940 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_198
timestamp 1644511149
transform 1 0 19320 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_205
timestamp 1644511149
transform 1 0 19964 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_218
timestamp 1644511149
transform 1 0 21160 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_225
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_236
timestamp 1644511149
transform 1 0 22816 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_244
timestamp 1644511149
transform 1 0 23552 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_254
timestamp 1644511149
transform 1 0 24472 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_265
timestamp 1644511149
transform 1 0 25484 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_274
timestamp 1644511149
transform 1 0 26312 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_289
timestamp 1644511149
transform 1 0 27692 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_296
timestamp 1644511149
transform 1 0 28336 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_308
timestamp 1644511149
transform 1 0 29440 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_320
timestamp 1644511149
transform 1 0 30544 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_332
timestamp 1644511149
transform 1 0 31648 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_349
timestamp 1644511149
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_361
timestamp 1644511149
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_373
timestamp 1644511149
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1644511149
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1644511149
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1644511149
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1644511149
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1644511149
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_61
timestamp 1644511149
transform 1 0 6716 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_78
timestamp 1644511149
transform 1 0 8280 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_96
timestamp 1644511149
transform 1 0 9936 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_106
timestamp 1644511149
transform 1 0 10856 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_114
timestamp 1644511149
transform 1 0 11592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_131
timestamp 1644511149
transform 1 0 13156 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1644511149
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_147
timestamp 1644511149
transform 1 0 14628 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_167
timestamp 1644511149
transform 1 0 16468 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_175
timestamp 1644511149
transform 1 0 17204 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_192
timestamp 1644511149
transform 1 0 18768 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_200
timestamp 1644511149
transform 1 0 19504 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_222
timestamp 1644511149
transform 1 0 21528 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_231
timestamp 1644511149
transform 1 0 22356 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_240
timestamp 1644511149
transform 1 0 23184 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_248
timestamp 1644511149
transform 1 0 23920 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_262
timestamp 1644511149
transform 1 0 25208 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_287
timestamp 1644511149
transform 1 0 27508 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_299
timestamp 1644511149
transform 1 0 28612 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1644511149
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_321
timestamp 1644511149
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_333
timestamp 1644511149
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_345
timestamp 1644511149
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1644511149
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1644511149
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_365
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_377
timestamp 1644511149
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_389
timestamp 1644511149
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_401
timestamp 1644511149
transform 1 0 37996 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1644511149
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1644511149
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1644511149
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1644511149
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1644511149
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_61
timestamp 1644511149
transform 1 0 6716 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_70
timestamp 1644511149
transform 1 0 7544 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_79
timestamp 1644511149
transform 1 0 8372 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_88
timestamp 1644511149
transform 1 0 9200 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_108
timestamp 1644511149
transform 1 0 11040 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_118
timestamp 1644511149
transform 1 0 11960 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_127
timestamp 1644511149
transform 1 0 12788 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_147
timestamp 1644511149
transform 1 0 14628 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_159
timestamp 1644511149
transform 1 0 15732 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1644511149
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_172
timestamp 1644511149
transform 1 0 16928 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_184
timestamp 1644511149
transform 1 0 18032 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_197
timestamp 1644511149
transform 1 0 19228 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_205
timestamp 1644511149
transform 1 0 19964 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_211
timestamp 1644511149
transform 1 0 20516 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_219
timestamp 1644511149
transform 1 0 21252 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1644511149
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_225
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_229
timestamp 1644511149
transform 1 0 22172 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_249
timestamp 1644511149
transform 1 0 24012 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_253
timestamp 1644511149
transform 1 0 24380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_260
timestamp 1644511149
transform 1 0 25024 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_274
timestamp 1644511149
transform 1 0 26312 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_293
timestamp 1644511149
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_305
timestamp 1644511149
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_317
timestamp 1644511149
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1644511149
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1644511149
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_349
timestamp 1644511149
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_361
timestamp 1644511149
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_373
timestamp 1644511149
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1644511149
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1644511149
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_405
timestamp 1644511149
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1644511149
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_61
timestamp 1644511149
transform 1 0 6716 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_80
timestamp 1644511149
transform 1 0 8464 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_88
timestamp 1644511149
transform 1 0 9200 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_99
timestamp 1644511149
transform 1 0 10212 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_111
timestamp 1644511149
transform 1 0 11316 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_125
timestamp 1644511149
transform 1 0 12604 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_134
timestamp 1644511149
transform 1 0 13432 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_153
timestamp 1644511149
transform 1 0 15180 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_173
timestamp 1644511149
transform 1 0 17020 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_179
timestamp 1644511149
transform 1 0 17572 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_192
timestamp 1644511149
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_209
timestamp 1644511149
transform 1 0 20332 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_225
timestamp 1644511149
transform 1 0 21804 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_238
timestamp 1644511149
transform 1 0 23000 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_247
timestamp 1644511149
transform 1 0 23828 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1644511149
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_253
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_265
timestamp 1644511149
transform 1 0 25484 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_273
timestamp 1644511149
transform 1 0 26220 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_285
timestamp 1644511149
transform 1 0 27324 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_297
timestamp 1644511149
transform 1 0 28428 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_305
timestamp 1644511149
transform 1 0 29164 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_321
timestamp 1644511149
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_333
timestamp 1644511149
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_345
timestamp 1644511149
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1644511149
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1644511149
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_377
timestamp 1644511149
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_389
timestamp 1644511149
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_401
timestamp 1644511149
transform 1 0 37996 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1644511149
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1644511149
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1644511149
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1644511149
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_75
timestamp 1644511149
transform 1 0 8004 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_97
timestamp 1644511149
transform 1 0 10028 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_109
timestamp 1644511149
transform 1 0 11132 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_119
timestamp 1644511149
transform 1 0 12052 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_139
timestamp 1644511149
transform 1 0 13892 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_161
timestamp 1644511149
transform 1 0 15916 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_177
timestamp 1644511149
transform 1 0 17388 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_184
timestamp 1644511149
transform 1 0 18032 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_188
timestamp 1644511149
transform 1 0 18400 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_192
timestamp 1644511149
transform 1 0 18768 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_196
timestamp 1644511149
transform 1 0 19136 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_200
timestamp 1644511149
transform 1 0 19504 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_204
timestamp 1644511149
transform 1 0 19872 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1644511149
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1644511149
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_225
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_240
timestamp 1644511149
transform 1 0 23184 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_260
timestamp 1644511149
transform 1 0 25024 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_267
timestamp 1644511149
transform 1 0 25668 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_274
timestamp 1644511149
transform 1 0 26312 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_293
timestamp 1644511149
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_305
timestamp 1644511149
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_317
timestamp 1644511149
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1644511149
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1644511149
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_337
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_349
timestamp 1644511149
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_361
timestamp 1644511149
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_373
timestamp 1644511149
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1644511149
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1644511149
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_405
timestamp 1644511149
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1644511149
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1644511149
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1644511149
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_93
timestamp 1644511149
transform 1 0 9660 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_111
timestamp 1644511149
transform 1 0 11316 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_119
timestamp 1644511149
transform 1 0 12052 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_129
timestamp 1644511149
transform 1 0 12972 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_136
timestamp 1644511149
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_144
timestamp 1644511149
transform 1 0 14352 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_151
timestamp 1644511149
transform 1 0 14996 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_155
timestamp 1644511149
transform 1 0 15364 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_172
timestamp 1644511149
transform 1 0 16928 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_180
timestamp 1644511149
transform 1 0 17664 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_185
timestamp 1644511149
transform 1 0 18124 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp 1644511149
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_197
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_210
timestamp 1644511149
transform 1 0 20424 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_218
timestamp 1644511149
transform 1 0 21160 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_233
timestamp 1644511149
transform 1 0 22540 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_239
timestamp 1644511149
transform 1 0 23092 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_243
timestamp 1644511149
transform 1 0 23460 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1644511149
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_253
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_280
timestamp 1644511149
transform 1 0 26864 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_292
timestamp 1644511149
transform 1 0 27968 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_304
timestamp 1644511149
transform 1 0 29072 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_321
timestamp 1644511149
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_333
timestamp 1644511149
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_345
timestamp 1644511149
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1644511149
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1644511149
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_377
timestamp 1644511149
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_389
timestamp 1644511149
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_401
timestamp 1644511149
transform 1 0 37996 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1644511149
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1644511149
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1644511149
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1644511149
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1644511149
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_93
timestamp 1644511149
transform 1 0 9660 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_97
timestamp 1644511149
transform 1 0 10028 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_102
timestamp 1644511149
transform 1 0 10488 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1644511149
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_121
timestamp 1644511149
transform 1 0 12236 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_129
timestamp 1644511149
transform 1 0 12972 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_138
timestamp 1644511149
transform 1 0 13800 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_158
timestamp 1644511149
transform 1 0 15640 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1644511149
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_176
timestamp 1644511149
transform 1 0 17296 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_185
timestamp 1644511149
transform 1 0 18124 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_193
timestamp 1644511149
transform 1 0 18860 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_202
timestamp 1644511149
transform 1 0 19688 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_213
timestamp 1644511149
transform 1 0 20700 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_220
timestamp 1644511149
transform 1 0 21344 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_237
timestamp 1644511149
transform 1 0 22908 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_255
timestamp 1644511149
transform 1 0 24564 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_271
timestamp 1644511149
transform 1 0 26036 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1644511149
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_281
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_293
timestamp 1644511149
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_305
timestamp 1644511149
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_317
timestamp 1644511149
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1644511149
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1644511149
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_349
timestamp 1644511149
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_361
timestamp 1644511149
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_373
timestamp 1644511149
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1644511149
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1644511149
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_393
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_405
timestamp 1644511149
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1644511149
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1644511149
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1644511149
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1644511149
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_97
timestamp 1644511149
transform 1 0 10028 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_106
timestamp 1644511149
transform 1 0 10856 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_113
timestamp 1644511149
transform 1 0 11500 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_125
timestamp 1644511149
transform 1 0 12604 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_137
timestamp 1644511149
transform 1 0 13708 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_146
timestamp 1644511149
transform 1 0 14536 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_159
timestamp 1644511149
transform 1 0 15732 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_163
timestamp 1644511149
transform 1 0 16100 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_174
timestamp 1644511149
transform 1 0 17112 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_183
timestamp 1644511149
transform 1 0 17940 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_191
timestamp 1644511149
transform 1 0 18676 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1644511149
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_209
timestamp 1644511149
transform 1 0 20332 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_218
timestamp 1644511149
transform 1 0 21160 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_234
timestamp 1644511149
transform 1 0 22632 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1644511149
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1644511149
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_258
timestamp 1644511149
transform 1 0 24840 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_266
timestamp 1644511149
transform 1 0 25576 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_273
timestamp 1644511149
transform 1 0 26220 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_281
timestamp 1644511149
transform 1 0 26956 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_290
timestamp 1644511149
transform 1 0 27784 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_302
timestamp 1644511149
transform 1 0 28888 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_309
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_317
timestamp 1644511149
transform 1 0 30268 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_324
timestamp 1644511149
transform 1 0 30912 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_331
timestamp 1644511149
transform 1 0 31556 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_337
timestamp 1644511149
transform 1 0 32108 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_341
timestamp 1644511149
transform 1 0 32476 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_353
timestamp 1644511149
transform 1 0 33580 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_361
timestamp 1644511149
transform 1 0 34316 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_365
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_377
timestamp 1644511149
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_389
timestamp 1644511149
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_401
timestamp 1644511149
transform 1 0 37996 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1644511149
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1644511149
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1644511149
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1644511149
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1644511149
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_89
timestamp 1644511149
transform 1 0 9292 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_106
timestamp 1644511149
transform 1 0 10856 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_121
timestamp 1644511149
transform 1 0 12236 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_125
timestamp 1644511149
transform 1 0 12604 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_134
timestamp 1644511149
transform 1 0 13432 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_142
timestamp 1644511149
transform 1 0 14168 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_150
timestamp 1644511149
transform 1 0 14904 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_155
timestamp 1644511149
transform 1 0 15364 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_164
timestamp 1644511149
transform 1 0 16192 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_178
timestamp 1644511149
transform 1 0 17480 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_186
timestamp 1644511149
transform 1 0 18216 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_190
timestamp 1644511149
transform 1 0 18584 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_201
timestamp 1644511149
transform 1 0 19596 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1644511149
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1644511149
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_228
timestamp 1644511149
transform 1 0 22080 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_234
timestamp 1644511149
transform 1 0 22632 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_247
timestamp 1644511149
transform 1 0 23828 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_254
timestamp 1644511149
transform 1 0 24472 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_262
timestamp 1644511149
transform 1 0 25208 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_268
timestamp 1644511149
transform 1 0 25760 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_276
timestamp 1644511149
transform 1 0 26496 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_281
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_296
timestamp 1644511149
transform 1 0 28336 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_306
timestamp 1644511149
transform 1 0 29256 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_318
timestamp 1644511149
transform 1 0 30360 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_328
timestamp 1644511149
transform 1 0 31280 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_342
timestamp 1644511149
transform 1 0 32568 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_351
timestamp 1644511149
transform 1 0 33396 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_362
timestamp 1644511149
transform 1 0 34408 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_369
timestamp 1644511149
transform 1 0 35052 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_381
timestamp 1644511149
transform 1 0 36156 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_389
timestamp 1644511149
transform 1 0 36892 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_393
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_405
timestamp 1644511149
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1644511149
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1644511149
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_73
timestamp 1644511149
transform 1 0 7820 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_79
timestamp 1644511149
transform 1 0 8372 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_94
timestamp 1644511149
transform 1 0 9752 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_105
timestamp 1644511149
transform 1 0 10764 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_115
timestamp 1644511149
transform 1 0 11684 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_119
timestamp 1644511149
transform 1 0 12052 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_136
timestamp 1644511149
transform 1 0 13616 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_141
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_160
timestamp 1644511149
transform 1 0 15824 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_172
timestamp 1644511149
transform 1 0 16928 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_180
timestamp 1644511149
transform 1 0 17664 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1644511149
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1644511149
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_201
timestamp 1644511149
transform 1 0 19596 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_222
timestamp 1644511149
transform 1 0 21528 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_238
timestamp 1644511149
transform 1 0 23000 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_248
timestamp 1644511149
transform 1 0 23920 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_261
timestamp 1644511149
transform 1 0 25116 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_273
timestamp 1644511149
transform 1 0 26220 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_283
timestamp 1644511149
transform 1 0 27140 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_291
timestamp 1644511149
transform 1 0 27876 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_299
timestamp 1644511149
transform 1 0 28612 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1644511149
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_317
timestamp 1644511149
transform 1 0 30268 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_327
timestamp 1644511149
transform 1 0 31188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_338
timestamp 1644511149
transform 1 0 32200 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_342
timestamp 1644511149
transform 1 0 32568 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_351
timestamp 1644511149
transform 1 0 33396 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_358
timestamp 1644511149
transform 1 0 34040 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_30_372
timestamp 1644511149
transform 1 0 35328 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_384
timestamp 1644511149
transform 1 0 36432 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_396
timestamp 1644511149
transform 1 0 37536 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_404
timestamp 1644511149
transform 1 0 38272 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1644511149
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1644511149
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1644511149
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1644511149
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1644511149
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_89
timestamp 1644511149
transform 1 0 9292 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_97
timestamp 1644511149
transform 1 0 10028 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_104
timestamp 1644511149
transform 1 0 10672 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_117
timestamp 1644511149
transform 1 0 11868 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_128
timestamp 1644511149
transform 1 0 12880 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_138
timestamp 1644511149
transform 1 0 13800 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_146
timestamp 1644511149
transform 1 0 14536 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_150
timestamp 1644511149
transform 1 0 14904 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_160
timestamp 1644511149
transform 1 0 15824 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_169
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_188
timestamp 1644511149
transform 1 0 18400 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_192
timestamp 1644511149
transform 1 0 18768 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_200
timestamp 1644511149
transform 1 0 19504 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_211
timestamp 1644511149
transform 1 0 20516 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_219
timestamp 1644511149
transform 1 0 21252 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1644511149
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_239
timestamp 1644511149
transform 1 0 23092 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_247
timestamp 1644511149
transform 1 0 23828 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_259
timestamp 1644511149
transform 1 0 24932 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_265
timestamp 1644511149
transform 1 0 25484 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_274
timestamp 1644511149
transform 1 0 26312 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_31_281
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_291
timestamp 1644511149
transform 1 0 27876 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_295
timestamp 1644511149
transform 1 0 28244 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_303
timestamp 1644511149
transform 1 0 28980 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_315
timestamp 1644511149
transform 1 0 30084 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_326
timestamp 1644511149
transform 1 0 31096 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_334
timestamp 1644511149
transform 1 0 31832 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_340
timestamp 1644511149
transform 1 0 32384 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_352
timestamp 1644511149
transform 1 0 33488 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_363
timestamp 1644511149
transform 1 0 34500 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_372
timestamp 1644511149
transform 1 0 35328 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_384
timestamp 1644511149
transform 1 0 36432 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_393
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1644511149
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1644511149
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_71
timestamp 1644511149
transform 1 0 7636 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_80
timestamp 1644511149
transform 1 0 8464 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_98
timestamp 1644511149
transform 1 0 10120 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_110
timestamp 1644511149
transform 1 0 11224 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_118
timestamp 1644511149
transform 1 0 11960 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_127
timestamp 1644511149
transform 1 0 12788 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_131
timestamp 1644511149
transform 1 0 13156 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_136
timestamp 1644511149
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_141
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_160
timestamp 1644511149
transform 1 0 15824 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_174
timestamp 1644511149
transform 1 0 17112 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_192
timestamp 1644511149
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_201
timestamp 1644511149
transform 1 0 19596 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_212
timestamp 1644511149
transform 1 0 20608 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_228
timestamp 1644511149
transform 1 0 22080 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_239
timestamp 1644511149
transform 1 0 23092 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_243
timestamp 1644511149
transform 1 0 23460 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_248
timestamp 1644511149
transform 1 0 23920 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_261
timestamp 1644511149
transform 1 0 25116 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_269
timestamp 1644511149
transform 1 0 25852 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_276
timestamp 1644511149
transform 1 0 26496 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_284
timestamp 1644511149
transform 1 0 27232 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_292
timestamp 1644511149
transform 1 0 27968 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_298
timestamp 1644511149
transform 1 0 28520 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_306
timestamp 1644511149
transform 1 0 29256 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_312
timestamp 1644511149
transform 1 0 29808 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_32_323
timestamp 1644511149
transform 1 0 30820 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_329
timestamp 1644511149
transform 1 0 31372 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_333
timestamp 1644511149
transform 1 0 31740 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_339
timestamp 1644511149
transform 1 0 32292 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_346
timestamp 1644511149
transform 1 0 32936 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_358
timestamp 1644511149
transform 1 0 34040 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_365
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_375
timestamp 1644511149
transform 1 0 35604 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_387
timestamp 1644511149
transform 1 0 36708 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_399
timestamp 1644511149
transform 1 0 37812 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1644511149
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1644511149
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1644511149
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1644511149
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_76
timestamp 1644511149
transform 1 0 8096 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_87
timestamp 1644511149
transform 1 0 9108 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_95
timestamp 1644511149
transform 1 0 9844 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_102
timestamp 1644511149
transform 1 0 10488 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1644511149
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_127
timestamp 1644511149
transform 1 0 12788 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_137
timestamp 1644511149
transform 1 0 13708 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_145
timestamp 1644511149
transform 1 0 14444 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_158
timestamp 1644511149
transform 1 0 15640 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1644511149
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_180
timestamp 1644511149
transform 1 0 17664 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_189
timestamp 1644511149
transform 1 0 18492 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_198
timestamp 1644511149
transform 1 0 19320 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_204
timestamp 1644511149
transform 1 0 19872 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1644511149
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1644511149
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_233
timestamp 1644511149
transform 1 0 22540 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_240
timestamp 1644511149
transform 1 0 23184 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_254
timestamp 1644511149
transform 1 0 24472 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_262
timestamp 1644511149
transform 1 0 25208 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_266
timestamp 1644511149
transform 1 0 25576 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_272
timestamp 1644511149
transform 1 0 26128 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_281
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_290
timestamp 1644511149
transform 1 0 27784 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_298
timestamp 1644511149
transform 1 0 28520 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_310
timestamp 1644511149
transform 1 0 29624 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_318
timestamp 1644511149
transform 1 0 30360 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_326
timestamp 1644511149
transform 1 0 31096 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_332
timestamp 1644511149
transform 1 0 31648 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_344
timestamp 1644511149
transform 1 0 32752 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_356
timestamp 1644511149
transform 1 0 33856 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_363
timestamp 1644511149
transform 1 0 34500 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_377
timestamp 1644511149
transform 1 0 35788 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_386
timestamp 1644511149
transform 1 0 36616 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_405
timestamp 1644511149
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_73
timestamp 1644511149
transform 1 0 7820 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_80
timestamp 1644511149
transform 1 0 8464 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_89
timestamp 1644511149
transform 1 0 9292 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_94
timestamp 1644511149
transform 1 0 9752 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_106
timestamp 1644511149
transform 1 0 10856 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_128
timestamp 1644511149
transform 1 0 12880 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_136
timestamp 1644511149
transform 1 0 13616 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_141
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_161
timestamp 1644511149
transform 1 0 15916 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_172
timestamp 1644511149
transform 1 0 16928 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_192
timestamp 1644511149
transform 1 0 18768 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_200
timestamp 1644511149
transform 1 0 19504 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_216
timestamp 1644511149
transform 1 0 20976 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_224
timestamp 1644511149
transform 1 0 21712 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_235
timestamp 1644511149
transform 1 0 22724 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_247
timestamp 1644511149
transform 1 0 23828 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1644511149
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_253
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_267
timestamp 1644511149
transform 1 0 25668 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_271
timestamp 1644511149
transform 1 0 26036 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_276
timestamp 1644511149
transform 1 0 26496 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_288
timestamp 1644511149
transform 1 0 27600 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_292
timestamp 1644511149
transform 1 0 27968 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_297
timestamp 1644511149
transform 1 0 28428 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_304
timestamp 1644511149
transform 1 0 29072 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_316
timestamp 1644511149
transform 1 0 30176 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_327
timestamp 1644511149
transform 1 0 31188 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_336
timestamp 1644511149
transform 1 0 32016 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_345
timestamp 1644511149
transform 1 0 32844 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_354
timestamp 1644511149
transform 1 0 33672 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_362
timestamp 1644511149
transform 1 0 34408 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_369
timestamp 1644511149
transform 1 0 35052 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_380
timestamp 1644511149
transform 1 0 36064 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_391
timestamp 1644511149
transform 1 0 37076 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_399
timestamp 1644511149
transform 1 0 37812 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1644511149
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1644511149
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1644511149
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1644511149
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1644511149
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_65
timestamp 1644511149
transform 1 0 7084 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_83
timestamp 1644511149
transform 1 0 8740 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_97
timestamp 1644511149
transform 1 0 10028 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1644511149
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1644511149
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_117
timestamp 1644511149
transform 1 0 11868 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_125
timestamp 1644511149
transform 1 0 12604 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_145
timestamp 1644511149
transform 1 0 14444 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_153
timestamp 1644511149
transform 1 0 15180 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_157
timestamp 1644511149
transform 1 0 15548 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_164
timestamp 1644511149
transform 1 0 16192 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_173
timestamp 1644511149
transform 1 0 17020 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_186
timestamp 1644511149
transform 1 0 18216 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_202
timestamp 1644511149
transform 1 0 19688 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_209
timestamp 1644511149
transform 1 0 20332 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_213
timestamp 1644511149
transform 1 0 20700 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1644511149
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1644511149
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_225
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_237
timestamp 1644511149
transform 1 0 22908 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_246
timestamp 1644511149
transform 1 0 23736 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_253
timestamp 1644511149
transform 1 0 24380 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_264
timestamp 1644511149
transform 1 0 25392 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_275
timestamp 1644511149
transform 1 0 26404 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1644511149
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_285
timestamp 1644511149
transform 1 0 27324 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_292
timestamp 1644511149
transform 1 0 27968 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_304
timestamp 1644511149
transform 1 0 29072 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_312
timestamp 1644511149
transform 1 0 29808 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_320
timestamp 1644511149
transform 1 0 30544 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_327
timestamp 1644511149
transform 1 0 31188 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1644511149
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_340
timestamp 1644511149
transform 1 0 32384 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_352
timestamp 1644511149
transform 1 0 33488 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_359
timestamp 1644511149
transform 1 0 34132 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_368
timestamp 1644511149
transform 1 0 34960 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_374
timestamp 1644511149
transform 1 0 35512 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1644511149
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1644511149
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_400
timestamp 1644511149
transform 1 0 37904 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_406
timestamp 1644511149
transform 1 0 38456 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_7
timestamp 1644511149
transform 1 0 1748 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_19
timestamp 1644511149
transform 1 0 2852 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_65
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1644511149
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1644511149
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_89
timestamp 1644511149
transform 1 0 9292 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_97
timestamp 1644511149
transform 1 0 10028 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_105
timestamp 1644511149
transform 1 0 10764 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_110
timestamp 1644511149
transform 1 0 11224 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_122
timestamp 1644511149
transform 1 0 12328 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_130
timestamp 1644511149
transform 1 0 13064 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_136
timestamp 1644511149
transform 1 0 13616 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_141
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_145
timestamp 1644511149
transform 1 0 14444 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_152
timestamp 1644511149
transform 1 0 15088 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_159
timestamp 1644511149
transform 1 0 15732 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_173
timestamp 1644511149
transform 1 0 17020 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_184
timestamp 1644511149
transform 1 0 18032 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_188
timestamp 1644511149
transform 1 0 18400 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_192
timestamp 1644511149
transform 1 0 18768 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_202
timestamp 1644511149
transform 1 0 19688 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_209
timestamp 1644511149
transform 1 0 20332 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_216
timestamp 1644511149
transform 1 0 20976 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_220
timestamp 1644511149
transform 1 0 21344 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_226
timestamp 1644511149
transform 1 0 21896 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_240
timestamp 1644511149
transform 1 0 23184 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_248
timestamp 1644511149
transform 1 0 23920 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_265
timestamp 1644511149
transform 1 0 25484 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_271
timestamp 1644511149
transform 1 0 26036 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_275
timestamp 1644511149
transform 1 0 26404 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_279
timestamp 1644511149
transform 1 0 26772 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_284
timestamp 1644511149
transform 1 0 27232 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_290
timestamp 1644511149
transform 1 0 27784 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_298
timestamp 1644511149
transform 1 0 28520 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_306
timestamp 1644511149
transform 1 0 29256 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_312
timestamp 1644511149
transform 1 0 29808 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_323
timestamp 1644511149
transform 1 0 30820 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_330
timestamp 1644511149
transform 1 0 31464 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_338
timestamp 1644511149
transform 1 0 32200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_343
timestamp 1644511149
transform 1 0 32660 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_347
timestamp 1644511149
transform 1 0 33028 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_354
timestamp 1644511149
transform 1 0 33672 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_362
timestamp 1644511149
transform 1 0 34408 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_369
timestamp 1644511149
transform 1 0 35052 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_376
timestamp 1644511149
transform 1 0 35696 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_388
timestamp 1644511149
transform 1 0 36800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_403
timestamp 1644511149
transform 1 0 38180 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1644511149
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1644511149
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1644511149
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1644511149
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_88
timestamp 1644511149
transform 1 0 9200 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_98
timestamp 1644511149
transform 1 0 10120 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1644511149
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1644511149
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_113
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_117
timestamp 1644511149
transform 1 0 11868 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_123
timestamp 1644511149
transform 1 0 12420 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_131
timestamp 1644511149
transform 1 0 13156 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_139
timestamp 1644511149
transform 1 0 13892 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_144
timestamp 1644511149
transform 1 0 14352 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_152
timestamp 1644511149
transform 1 0 15088 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_156
timestamp 1644511149
transform 1 0 15456 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1644511149
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1644511149
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_175
timestamp 1644511149
transform 1 0 17204 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_182
timestamp 1644511149
transform 1 0 17848 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_189
timestamp 1644511149
transform 1 0 18492 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_37_200
timestamp 1644511149
transform 1 0 19504 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_220
timestamp 1644511149
transform 1 0 21344 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_236
timestamp 1644511149
transform 1 0 22816 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_240
timestamp 1644511149
transform 1 0 23184 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_248
timestamp 1644511149
transform 1 0 23920 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_259
timestamp 1644511149
transform 1 0 24932 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_37_270
timestamp 1644511149
transform 1 0 25944 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_278
timestamp 1644511149
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_289
timestamp 1644511149
transform 1 0 27692 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_295
timestamp 1644511149
transform 1 0 28244 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_301
timestamp 1644511149
transform 1 0 28796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_308
timestamp 1644511149
transform 1 0 29440 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_315
timestamp 1644511149
transform 1 0 30084 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_319
timestamp 1644511149
transform 1 0 30452 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_323
timestamp 1644511149
transform 1 0 30820 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_331
timestamp 1644511149
transform 1 0 31556 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1644511149
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_340
timestamp 1644511149
transform 1 0 32384 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_349
timestamp 1644511149
transform 1 0 33212 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_358
timestamp 1644511149
transform 1 0 34040 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_366
timestamp 1644511149
transform 1 0 34776 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_376
timestamp 1644511149
transform 1 0 35696 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1644511149
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1644511149
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_393
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_405
timestamp 1644511149
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1644511149
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1644511149
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_61
timestamp 1644511149
transform 1 0 6716 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_80
timestamp 1644511149
transform 1 0 8464 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_92
timestamp 1644511149
transform 1 0 9568 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_104
timestamp 1644511149
transform 1 0 10672 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_115
timestamp 1644511149
transform 1 0 11684 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_38_131
timestamp 1644511149
transform 1 0 13156 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1644511149
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_158
timestamp 1644511149
transform 1 0 15640 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_166
timestamp 1644511149
transform 1 0 16376 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_174
timestamp 1644511149
transform 1 0 17112 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_182
timestamp 1644511149
transform 1 0 17848 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_188
timestamp 1644511149
transform 1 0 18400 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_192
timestamp 1644511149
transform 1 0 18768 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_202
timestamp 1644511149
transform 1 0 19688 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_223
timestamp 1644511149
transform 1 0 21620 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_239
timestamp 1644511149
transform 1 0 23092 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_247
timestamp 1644511149
transform 1 0 23828 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1644511149
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_260
timestamp 1644511149
transform 1 0 25024 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_267
timestamp 1644511149
transform 1 0 25668 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_275
timestamp 1644511149
transform 1 0 26404 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_282
timestamp 1644511149
transform 1 0 27048 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_291
timestamp 1644511149
transform 1 0 27876 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1644511149
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1644511149
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_309
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_313
timestamp 1644511149
transform 1 0 29900 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_324
timestamp 1644511149
transform 1 0 30912 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_335
timestamp 1644511149
transform 1 0 31924 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_343
timestamp 1644511149
transform 1 0 32660 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_349
timestamp 1644511149
transform 1 0 33212 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1644511149
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1644511149
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_365
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_372
timestamp 1644511149
transform 1 0 35328 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_381
timestamp 1644511149
transform 1 0 36156 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_385
timestamp 1644511149
transform 1 0 36524 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_392
timestamp 1644511149
transform 1 0 37168 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_399
timestamp 1644511149
transform 1 0 37812 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1644511149
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1644511149
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1644511149
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1644511149
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_77
timestamp 1644511149
transform 1 0 8188 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_82
timestamp 1644511149
transform 1 0 8648 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_93
timestamp 1644511149
transform 1 0 9660 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_101
timestamp 1644511149
transform 1 0 10396 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_109
timestamp 1644511149
transform 1 0 11132 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_123
timestamp 1644511149
transform 1 0 12420 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_130
timestamp 1644511149
transform 1 0 13064 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_137
timestamp 1644511149
transform 1 0 13708 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_146
timestamp 1644511149
transform 1 0 14536 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_153
timestamp 1644511149
transform 1 0 15180 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_162
timestamp 1644511149
transform 1 0 16008 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_174
timestamp 1644511149
transform 1 0 17112 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_178
timestamp 1644511149
transform 1 0 17480 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_184
timestamp 1644511149
transform 1 0 18032 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_192
timestamp 1644511149
transform 1 0 18768 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_199
timestamp 1644511149
transform 1 0 19412 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_208
timestamp 1644511149
transform 1 0 20240 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_216
timestamp 1644511149
transform 1 0 20976 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_220
timestamp 1644511149
transform 1 0 21344 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_225
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_229
timestamp 1644511149
transform 1 0 22172 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_236
timestamp 1644511149
transform 1 0 22816 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_247
timestamp 1644511149
transform 1 0 23828 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_254
timestamp 1644511149
transform 1 0 24472 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_39_270
timestamp 1644511149
transform 1 0 25944 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_278
timestamp 1644511149
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_281
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_287
timestamp 1644511149
transform 1 0 27508 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_294
timestamp 1644511149
transform 1 0 28152 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_305
timestamp 1644511149
transform 1 0 29164 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_313
timestamp 1644511149
transform 1 0 29900 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_331
timestamp 1644511149
transform 1 0 31556 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1644511149
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_337
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_343
timestamp 1644511149
transform 1 0 32660 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_350
timestamp 1644511149
transform 1 0 33304 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_358
timestamp 1644511149
transform 1 0 34040 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_368
timestamp 1644511149
transform 1 0 34960 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_378
timestamp 1644511149
transform 1 0 35880 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_386
timestamp 1644511149
transform 1 0 36616 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_39_400
timestamp 1644511149
transform 1 0 37904 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_406
timestamp 1644511149
transform 1 0 38456 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1644511149
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_109
timestamp 1644511149
transform 1 0 11132 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_119
timestamp 1644511149
transform 1 0 12052 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_130
timestamp 1644511149
transform 1 0 13064 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1644511149
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_146
timestamp 1644511149
transform 1 0 14536 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_155
timestamp 1644511149
transform 1 0 15364 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_164
timestamp 1644511149
transform 1 0 16192 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_173
timestamp 1644511149
transform 1 0 17020 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_177
timestamp 1644511149
transform 1 0 17388 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_183
timestamp 1644511149
transform 1 0 17940 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_190
timestamp 1644511149
transform 1 0 18584 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_204
timestamp 1644511149
transform 1 0 19872 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_208
timestamp 1644511149
transform 1 0 20240 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_212
timestamp 1644511149
transform 1 0 20608 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_228
timestamp 1644511149
transform 1 0 22080 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_236
timestamp 1644511149
transform 1 0 22816 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1644511149
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1644511149
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_253
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_257
timestamp 1644511149
transform 1 0 24748 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_264
timestamp 1644511149
transform 1 0 25392 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_271
timestamp 1644511149
transform 1 0 26036 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_283
timestamp 1644511149
transform 1 0 27140 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_290
timestamp 1644511149
transform 1 0 27784 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_298
timestamp 1644511149
transform 1 0 28520 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_303
timestamp 1644511149
transform 1 0 28980 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1644511149
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_314
timestamp 1644511149
transform 1 0 29992 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_321
timestamp 1644511149
transform 1 0 30636 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_40_330
timestamp 1644511149
transform 1 0 31464 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_342
timestamp 1644511149
transform 1 0 32568 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_356
timestamp 1644511149
transform 1 0 33856 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_368
timestamp 1644511149
transform 1 0 34960 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_375
timestamp 1644511149
transform 1 0 35604 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_388
timestamp 1644511149
transform 1 0 36800 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_399
timestamp 1644511149
transform 1 0 37812 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1644511149
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1644511149
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1644511149
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_81
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_93
timestamp 1644511149
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1644511149
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1644511149
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_125
timestamp 1644511149
transform 1 0 12604 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_138
timestamp 1644511149
transform 1 0 13800 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_147
timestamp 1644511149
transform 1 0 14628 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_156
timestamp 1644511149
transform 1 0 15456 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_160
timestamp 1644511149
transform 1 0 15824 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_164
timestamp 1644511149
transform 1 0 16192 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_183
timestamp 1644511149
transform 1 0 17940 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_199
timestamp 1644511149
transform 1 0 19412 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_206
timestamp 1644511149
transform 1 0 20056 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_213
timestamp 1644511149
transform 1 0 20700 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_220
timestamp 1644511149
transform 1 0 21344 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_237
timestamp 1644511149
transform 1 0 22908 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_241
timestamp 1644511149
transform 1 0 23276 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_246
timestamp 1644511149
transform 1 0 23736 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_250
timestamp 1644511149
transform 1 0 24104 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_256
timestamp 1644511149
transform 1 0 24656 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_268
timestamp 1644511149
transform 1 0 25760 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_276
timestamp 1644511149
transform 1 0 26496 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_286
timestamp 1644511149
transform 1 0 27416 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_314
timestamp 1644511149
transform 1 0 29992 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_328
timestamp 1644511149
transform 1 0 31280 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_340
timestamp 1644511149
transform 1 0 32384 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_347
timestamp 1644511149
transform 1 0 33028 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_353
timestamp 1644511149
transform 1 0 33580 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_362
timestamp 1644511149
transform 1 0 34408 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_371
timestamp 1644511149
transform 1 0 35236 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_377
timestamp 1644511149
transform 1 0 35788 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_383
timestamp 1644511149
transform 1 0 36340 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1644511149
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_399
timestamp 1644511149
transform 1 0 37812 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1644511149
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1644511149
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1644511149
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1644511149
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1644511149
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_97
timestamp 1644511149
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_109
timestamp 1644511149
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_121
timestamp 1644511149
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_136
timestamp 1644511149
transform 1 0 13616 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_144
timestamp 1644511149
transform 1 0 14352 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_155
timestamp 1644511149
transform 1 0 15364 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_162
timestamp 1644511149
transform 1 0 16008 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_178
timestamp 1644511149
transform 1 0 17480 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_186
timestamp 1644511149
transform 1 0 18216 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_191
timestamp 1644511149
transform 1 0 18676 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1644511149
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_197
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_213
timestamp 1644511149
transform 1 0 20700 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_220
timestamp 1644511149
transform 1 0 21344 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_42_237
timestamp 1644511149
transform 1 0 22908 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_243
timestamp 1644511149
transform 1 0 23460 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_248
timestamp 1644511149
transform 1 0 23920 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_263
timestamp 1644511149
transform 1 0 25300 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_271
timestamp 1644511149
transform 1 0 26036 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_279
timestamp 1644511149
transform 1 0 26772 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_285
timestamp 1644511149
transform 1 0 27324 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_291
timestamp 1644511149
transform 1 0 27876 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_299
timestamp 1644511149
transform 1 0 28612 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1644511149
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_316
timestamp 1644511149
transform 1 0 30176 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_325
timestamp 1644511149
transform 1 0 31004 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_332
timestamp 1644511149
transform 1 0 31648 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_340
timestamp 1644511149
transform 1 0 32384 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_344
timestamp 1644511149
transform 1 0 32752 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_360
timestamp 1644511149
transform 1 0 34224 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_373
timestamp 1644511149
transform 1 0 35420 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_382
timestamp 1644511149
transform 1 0 36248 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_390
timestamp 1644511149
transform 1 0 36984 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_42_400
timestamp 1644511149
transform 1 0 37904 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_406
timestamp 1644511149
transform 1 0 38456 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1644511149
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1644511149
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1644511149
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1644511149
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_93
timestamp 1644511149
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1644511149
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_125
timestamp 1644511149
transform 1 0 12604 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_134
timestamp 1644511149
transform 1 0 13432 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_141
timestamp 1644511149
transform 1 0 14076 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_148
timestamp 1644511149
transform 1 0 14720 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_164
timestamp 1644511149
transform 1 0 16192 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_181
timestamp 1644511149
transform 1 0 17756 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_189
timestamp 1644511149
transform 1 0 18492 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_197
timestamp 1644511149
transform 1 0 19228 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_201
timestamp 1644511149
transform 1 0 19596 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_209
timestamp 1644511149
transform 1 0 20332 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_216
timestamp 1644511149
transform 1 0 20976 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_43_225
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_235
timestamp 1644511149
transform 1 0 22724 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_243
timestamp 1644511149
transform 1 0 23460 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_252
timestamp 1644511149
transform 1 0 24288 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_263
timestamp 1644511149
transform 1 0 25300 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_275
timestamp 1644511149
transform 1 0 26404 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1644511149
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_281
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_285
timestamp 1644511149
transform 1 0 27324 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_290
timestamp 1644511149
transform 1 0 27784 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_302
timestamp 1644511149
transform 1 0 28888 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_306
timestamp 1644511149
transform 1 0 29256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_312
timestamp 1644511149
transform 1 0 29808 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_322
timestamp 1644511149
transform 1 0 30728 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1644511149
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1644511149
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_337
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_346
timestamp 1644511149
transform 1 0 32936 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_357
timestamp 1644511149
transform 1 0 33948 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_365
timestamp 1644511149
transform 1 0 34684 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_369
timestamp 1644511149
transform 1 0 35052 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_374
timestamp 1644511149
transform 1 0 35512 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_382
timestamp 1644511149
transform 1 0 36248 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_390
timestamp 1644511149
transform 1 0 36984 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_400
timestamp 1644511149
transform 1 0 37904 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_406
timestamp 1644511149
transform 1 0 38456 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1644511149
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1644511149
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_97
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_109
timestamp 1644511149
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_121
timestamp 1644511149
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1644511149
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1644511149
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_155
timestamp 1644511149
transform 1 0 15364 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_171
timestamp 1644511149
transform 1 0 16836 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_179
timestamp 1644511149
transform 1 0 17572 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_188
timestamp 1644511149
transform 1 0 18400 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_197
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_201
timestamp 1644511149
transform 1 0 19596 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_209
timestamp 1644511149
transform 1 0 20332 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_217
timestamp 1644511149
transform 1 0 21068 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_227
timestamp 1644511149
transform 1 0 21988 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_248
timestamp 1644511149
transform 1 0 23920 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_253
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_44_262
timestamp 1644511149
transform 1 0 25208 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_272
timestamp 1644511149
transform 1 0 26128 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_280
timestamp 1644511149
transform 1 0 26864 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_291
timestamp 1644511149
transform 1 0 27876 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_299
timestamp 1644511149
transform 1 0 28612 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1644511149
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_312
timestamp 1644511149
transform 1 0 29808 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_316
timestamp 1644511149
transform 1 0 30176 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_324
timestamp 1644511149
transform 1 0 30912 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_332
timestamp 1644511149
transform 1 0 31648 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_337
timestamp 1644511149
transform 1 0 32108 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_348
timestamp 1644511149
transform 1 0 33120 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_44_358
timestamp 1644511149
transform 1 0 34040 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_372
timestamp 1644511149
transform 1 0 35328 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_382
timestamp 1644511149
transform 1 0 36248 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_403
timestamp 1644511149
transform 1 0 38180 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1644511149
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1644511149
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1644511149
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1644511149
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1644511149
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_93
timestamp 1644511149
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1644511149
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1644511149
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_125
timestamp 1644511149
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_137
timestamp 1644511149
transform 1 0 13708 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_143
timestamp 1644511149
transform 1 0 14260 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_156
timestamp 1644511149
transform 1 0 15456 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_160
timestamp 1644511149
transform 1 0 15824 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_164
timestamp 1644511149
transform 1 0 16192 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_176
timestamp 1644511149
transform 1 0 17296 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_187
timestamp 1644511149
transform 1 0 18308 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_195
timestamp 1644511149
transform 1 0 19044 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_203
timestamp 1644511149
transform 1 0 19780 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_211
timestamp 1644511149
transform 1 0 20516 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_215
timestamp 1644511149
transform 1 0 20884 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_220
timestamp 1644511149
transform 1 0 21344 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_225
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_229
timestamp 1644511149
transform 1 0 22172 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_238
timestamp 1644511149
transform 1 0 23000 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_246
timestamp 1644511149
transform 1 0 23736 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_253
timestamp 1644511149
transform 1 0 24380 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_262
timestamp 1644511149
transform 1 0 25208 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_271
timestamp 1644511149
transform 1 0 26036 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1644511149
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_291
timestamp 1644511149
transform 1 0 27876 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_302
timestamp 1644511149
transform 1 0 28888 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_317
timestamp 1644511149
transform 1 0 30268 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1644511149
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1644511149
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_344
timestamp 1644511149
transform 1 0 32752 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_356
timestamp 1644511149
transform 1 0 33856 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_360
timestamp 1644511149
transform 1 0 34224 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_369
timestamp 1644511149
transform 1 0 35052 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_380
timestamp 1644511149
transform 1 0 36064 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_387
timestamp 1644511149
transform 1 0 36708 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1644511149
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_400
timestamp 1644511149
transform 1 0 37904 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_406
timestamp 1644511149
transform 1 0 38456 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_65
timestamp 1644511149
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1644511149
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1644511149
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_97
timestamp 1644511149
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_109
timestamp 1644511149
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_121
timestamp 1644511149
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1644511149
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1644511149
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_157
timestamp 1644511149
transform 1 0 15548 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_163
timestamp 1644511149
transform 1 0 16100 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_168
timestamp 1644511149
transform 1 0 16560 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_176
timestamp 1644511149
transform 1 0 17296 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_180
timestamp 1644511149
transform 1 0 17664 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_188
timestamp 1644511149
transform 1 0 18400 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_201
timestamp 1644511149
transform 1 0 19596 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_211
timestamp 1644511149
transform 1 0 20516 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_215
timestamp 1644511149
transform 1 0 20884 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_220
timestamp 1644511149
transform 1 0 21344 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_224
timestamp 1644511149
transform 1 0 21712 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_230
timestamp 1644511149
transform 1 0 22264 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_46_243
timestamp 1644511149
transform 1 0 23460 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1644511149
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_253
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_263
timestamp 1644511149
transform 1 0 25300 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_271
timestamp 1644511149
transform 1 0 26036 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_279
timestamp 1644511149
transform 1 0 26772 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_290
timestamp 1644511149
transform 1 0 27784 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_299
timestamp 1644511149
transform 1 0 28612 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1644511149
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_313
timestamp 1644511149
transform 1 0 29900 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_320
timestamp 1644511149
transform 1 0 30544 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_327
timestamp 1644511149
transform 1 0 31188 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_46_342
timestamp 1644511149
transform 1 0 32568 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_350
timestamp 1644511149
transform 1 0 33304 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_360
timestamp 1644511149
transform 1 0 34224 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_369
timestamp 1644511149
transform 1 0 35052 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_376
timestamp 1644511149
transform 1 0 35696 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_387
timestamp 1644511149
transform 1 0 36708 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_394
timestamp 1644511149
transform 1 0 37352 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_401
timestamp 1644511149
transform 1 0 37996 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1644511149
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1644511149
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1644511149
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_93
timestamp 1644511149
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1644511149
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1644511149
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_125
timestamp 1644511149
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_137
timestamp 1644511149
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1644511149
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1644511149
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_47_169
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_177
timestamp 1644511149
transform 1 0 17388 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_185
timestamp 1644511149
transform 1 0 18124 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_195
timestamp 1644511149
transform 1 0 19044 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_206
timestamp 1644511149
transform 1 0 20056 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_218
timestamp 1644511149
transform 1 0 21160 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_228
timestamp 1644511149
transform 1 0 22080 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_236
timestamp 1644511149
transform 1 0 22816 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_244
timestamp 1644511149
transform 1 0 23552 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_252
timestamp 1644511149
transform 1 0 24288 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_260
timestamp 1644511149
transform 1 0 25024 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1644511149
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1644511149
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_281
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_289
timestamp 1644511149
transform 1 0 27692 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_299
timestamp 1644511149
transform 1 0 28612 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_308
timestamp 1644511149
transform 1 0 29440 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_316
timestamp 1644511149
transform 1 0 30176 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_322
timestamp 1644511149
transform 1 0 30728 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_330
timestamp 1644511149
transform 1 0 31464 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_47_344
timestamp 1644511149
transform 1 0 32752 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_352
timestamp 1644511149
transform 1 0 33488 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_357
timestamp 1644511149
transform 1 0 33948 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_364
timestamp 1644511149
transform 1 0 34592 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_371
timestamp 1644511149
transform 1 0 35236 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_377
timestamp 1644511149
transform 1 0 35788 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_381
timestamp 1644511149
transform 1 0 36156 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_388
timestamp 1644511149
transform 1 0 36800 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_393
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_399
timestamp 1644511149
transform 1 0 37812 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1644511149
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_109
timestamp 1644511149
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_121
timestamp 1644511149
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1644511149
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1644511149
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_141
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_153
timestamp 1644511149
transform 1 0 15180 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_159
timestamp 1644511149
transform 1 0 15732 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_168
timestamp 1644511149
transform 1 0 16560 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_181
timestamp 1644511149
transform 1 0 17756 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_192
timestamp 1644511149
transform 1 0 18768 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_210
timestamp 1644511149
transform 1 0 20424 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_221
timestamp 1644511149
transform 1 0 21436 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_228
timestamp 1644511149
transform 1 0 22080 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_234
timestamp 1644511149
transform 1 0 22632 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_239
timestamp 1644511149
transform 1 0 23092 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_248
timestamp 1644511149
transform 1 0 23920 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_253
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_261
timestamp 1644511149
transform 1 0 25116 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_269
timestamp 1644511149
transform 1 0 25852 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_276
timestamp 1644511149
transform 1 0 26496 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_282
timestamp 1644511149
transform 1 0 27048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_290
timestamp 1644511149
transform 1 0 27784 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_304
timestamp 1644511149
transform 1 0 29072 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_309
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_319
timestamp 1644511149
transform 1 0 30452 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_326
timestamp 1644511149
transform 1 0 31096 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_334
timestamp 1644511149
transform 1 0 31832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_339
timestamp 1644511149
transform 1 0 32292 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_346
timestamp 1644511149
transform 1 0 32936 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_353
timestamp 1644511149
transform 1 0 33580 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_360
timestamp 1644511149
transform 1 0 34224 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_369
timestamp 1644511149
transform 1 0 35052 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_48_382
timestamp 1644511149
transform 1 0 36248 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_394
timestamp 1644511149
transform 1 0 37352 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_403
timestamp 1644511149
transform 1 0 38180 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1644511149
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1644511149
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1644511149
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1644511149
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_93
timestamp 1644511149
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1644511149
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_125
timestamp 1644511149
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_137
timestamp 1644511149
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_149
timestamp 1644511149
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_164
timestamp 1644511149
transform 1 0 16192 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_173
timestamp 1644511149
transform 1 0 17020 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_183
timestamp 1644511149
transform 1 0 17940 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_190
timestamp 1644511149
transform 1 0 18584 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_198
timestamp 1644511149
transform 1 0 19320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_209
timestamp 1644511149
transform 1 0 20332 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_216
timestamp 1644511149
transform 1 0 20976 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_225
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_233
timestamp 1644511149
transform 1 0 22540 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_240
timestamp 1644511149
transform 1 0 23184 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_244
timestamp 1644511149
transform 1 0 23552 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_252
timestamp 1644511149
transform 1 0 24288 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_262
timestamp 1644511149
transform 1 0 25208 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_49_274
timestamp 1644511149
transform 1 0 26312 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_281
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_285
timestamp 1644511149
transform 1 0 27324 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_294
timestamp 1644511149
transform 1 0 28152 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_303
timestamp 1644511149
transform 1 0 28980 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_307
timestamp 1644511149
transform 1 0 29348 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_315
timestamp 1644511149
transform 1 0 30084 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_322
timestamp 1644511149
transform 1 0 30728 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_330
timestamp 1644511149
transform 1 0 31464 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_342
timestamp 1644511149
transform 1 0 32568 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_350
timestamp 1644511149
transform 1 0 33304 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_361
timestamp 1644511149
transform 1 0 34316 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_370
timestamp 1644511149
transform 1 0 35144 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_379
timestamp 1644511149
transform 1 0 35972 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_383
timestamp 1644511149
transform 1 0 36340 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_388
timestamp 1644511149
transform 1 0 36800 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_401
timestamp 1644511149
transform 1 0 37996 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1644511149
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1644511149
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1644511149
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_97
timestamp 1644511149
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_109
timestamp 1644511149
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_121
timestamp 1644511149
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1644511149
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1644511149
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_153
timestamp 1644511149
transform 1 0 15180 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_162
timestamp 1644511149
transform 1 0 16008 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_176
timestamp 1644511149
transform 1 0 17296 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_182
timestamp 1644511149
transform 1 0 17848 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_188
timestamp 1644511149
transform 1 0 18400 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_50_197
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_50_208
timestamp 1644511149
transform 1 0 20240 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_216
timestamp 1644511149
transform 1 0 20976 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_221
timestamp 1644511149
transform 1 0 21436 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_229
timestamp 1644511149
transform 1 0 22172 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_238
timestamp 1644511149
transform 1 0 23000 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_247
timestamp 1644511149
transform 1 0 23828 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1644511149
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_257
timestamp 1644511149
transform 1 0 24748 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_268
timestamp 1644511149
transform 1 0 25760 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_277
timestamp 1644511149
transform 1 0 26588 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_285
timestamp 1644511149
transform 1 0 27324 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_300
timestamp 1644511149
transform 1 0 28704 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_309
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_317
timestamp 1644511149
transform 1 0 30268 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_321
timestamp 1644511149
transform 1 0 30636 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_326
timestamp 1644511149
transform 1 0 31096 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_344
timestamp 1644511149
transform 1 0 32752 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_355
timestamp 1644511149
transform 1 0 33764 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1644511149
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_368
timestamp 1644511149
transform 1 0 34960 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_375
timestamp 1644511149
transform 1 0 35604 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_379
timestamp 1644511149
transform 1 0 35972 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_384
timestamp 1644511149
transform 1 0 36432 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_396
timestamp 1644511149
transform 1 0 37536 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_404
timestamp 1644511149
transform 1 0 38272 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1644511149
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1644511149
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1644511149
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1644511149
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1644511149
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1644511149
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1644511149
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_125
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_137
timestamp 1644511149
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_149
timestamp 1644511149
transform 1 0 14812 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_164
timestamp 1644511149
transform 1 0 16192 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_190
timestamp 1644511149
transform 1 0 18584 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_201
timestamp 1644511149
transform 1 0 19596 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_209
timestamp 1644511149
transform 1 0 20332 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_216
timestamp 1644511149
transform 1 0 20976 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_230
timestamp 1644511149
transform 1 0 22264 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_239
timestamp 1644511149
transform 1 0 23092 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_247
timestamp 1644511149
transform 1 0 23828 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_251
timestamp 1644511149
transform 1 0 24196 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_257
timestamp 1644511149
transform 1 0 24748 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_274
timestamp 1644511149
transform 1 0 26312 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_281
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_285
timestamp 1644511149
transform 1 0 27324 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_294
timestamp 1644511149
transform 1 0 28152 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_51_304
timestamp 1644511149
transform 1 0 29072 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_312
timestamp 1644511149
transform 1 0 29808 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_324
timestamp 1644511149
transform 1 0 30912 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_332
timestamp 1644511149
transform 1 0 31648 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_341
timestamp 1644511149
transform 1 0 32476 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_348
timestamp 1644511149
transform 1 0 33120 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_356
timestamp 1644511149
transform 1 0 33856 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_363
timestamp 1644511149
transform 1 0 34500 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_371
timestamp 1644511149
transform 1 0 35236 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_379
timestamp 1644511149
transform 1 0 35972 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_387
timestamp 1644511149
transform 1 0 36708 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1644511149
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_400
timestamp 1644511149
transform 1 0 37904 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_406
timestamp 1644511149
transform 1 0 38456 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1644511149
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1644511149
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_121
timestamp 1644511149
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1644511149
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_161
timestamp 1644511149
transform 1 0 15916 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_174
timestamp 1644511149
transform 1 0 17112 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_52_190
timestamp 1644511149
transform 1 0 18584 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_52_203
timestamp 1644511149
transform 1 0 19780 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_214
timestamp 1644511149
transform 1 0 20792 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_218
timestamp 1644511149
transform 1 0 21160 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_225
timestamp 1644511149
transform 1 0 21804 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_232
timestamp 1644511149
transform 1 0 22448 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_236
timestamp 1644511149
transform 1 0 22816 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_244
timestamp 1644511149
transform 1 0 23552 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_52_253
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_52_265
timestamp 1644511149
transform 1 0 25484 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_274
timestamp 1644511149
transform 1 0 26312 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_285
timestamp 1644511149
transform 1 0 27324 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_291
timestamp 1644511149
transform 1 0 27876 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_296
timestamp 1644511149
transform 1 0 28336 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_304
timestamp 1644511149
transform 1 0 29072 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_313
timestamp 1644511149
transform 1 0 29900 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_322
timestamp 1644511149
transform 1 0 30728 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_335
timestamp 1644511149
transform 1 0 31924 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_344
timestamp 1644511149
transform 1 0 32752 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_350
timestamp 1644511149
transform 1 0 33304 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_354
timestamp 1644511149
transform 1 0 33672 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_362
timestamp 1644511149
transform 1 0 34408 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_365
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_372
timestamp 1644511149
transform 1 0 35328 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_383
timestamp 1644511149
transform 1 0 36340 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_395
timestamp 1644511149
transform 1 0 37444 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_15
timestamp 1644511149
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_27
timestamp 1644511149
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_39
timestamp 1644511149
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1644511149
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1644511149
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_93
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1644511149
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1644511149
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_125
timestamp 1644511149
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_137
timestamp 1644511149
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_149
timestamp 1644511149
transform 1 0 14812 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_155
timestamp 1644511149
transform 1 0 15364 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_164
timestamp 1644511149
transform 1 0 16192 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_169
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_178
timestamp 1644511149
transform 1 0 17480 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_182
timestamp 1644511149
transform 1 0 17848 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_188
timestamp 1644511149
transform 1 0 18400 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_198
timestamp 1644511149
transform 1 0 19320 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_212
timestamp 1644511149
transform 1 0 20608 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_219
timestamp 1644511149
transform 1 0 21252 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1644511149
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_232
timestamp 1644511149
transform 1 0 22448 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_243
timestamp 1644511149
transform 1 0 23460 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_250
timestamp 1644511149
transform 1 0 24104 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_257
timestamp 1644511149
transform 1 0 24748 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_265
timestamp 1644511149
transform 1 0 25484 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_276
timestamp 1644511149
transform 1 0 26496 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_289
timestamp 1644511149
transform 1 0 27692 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_300
timestamp 1644511149
transform 1 0 28704 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_307
timestamp 1644511149
transform 1 0 29348 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_316
timestamp 1644511149
transform 1 0 30176 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1644511149
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1644511149
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_337
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_341
timestamp 1644511149
transform 1 0 32476 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_349
timestamp 1644511149
transform 1 0 33212 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_356
timestamp 1644511149
transform 1 0 33856 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_360
timestamp 1644511149
transform 1 0 34224 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_368
timestamp 1644511149
transform 1 0 34960 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_379
timestamp 1644511149
transform 1 0 35972 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1644511149
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_393
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_405
timestamp 1644511149
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_15
timestamp 1644511149
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1644511149
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1644511149
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1644511149
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1644511149
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1644511149
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_121
timestamp 1644511149
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1644511149
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1644511149
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_141
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_153
timestamp 1644511149
transform 1 0 15180 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_157
timestamp 1644511149
transform 1 0 15548 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_166
timestamp 1644511149
transform 1 0 16376 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_174
timestamp 1644511149
transform 1 0 17112 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_182
timestamp 1644511149
transform 1 0 17848 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_192
timestamp 1644511149
transform 1 0 18768 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_204
timestamp 1644511149
transform 1 0 19872 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_54_218
timestamp 1644511149
transform 1 0 21160 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_54_231
timestamp 1644511149
transform 1 0 22356 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_248
timestamp 1644511149
transform 1 0 23920 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_260
timestamp 1644511149
transform 1 0 25024 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_264
timestamp 1644511149
transform 1 0 25392 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_274
timestamp 1644511149
transform 1 0 26312 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_282
timestamp 1644511149
transform 1 0 27048 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_286
timestamp 1644511149
transform 1 0 27416 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_291
timestamp 1644511149
transform 1 0 27876 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_300
timestamp 1644511149
transform 1 0 28704 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_319
timestamp 1644511149
transform 1 0 30452 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_323
timestamp 1644511149
transform 1 0 30820 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_332
timestamp 1644511149
transform 1 0 31648 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_343
timestamp 1644511149
transform 1 0 32660 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_347
timestamp 1644511149
transform 1 0 33028 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_353
timestamp 1644511149
transform 1 0 33580 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_360
timestamp 1644511149
transform 1 0 34224 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_368
timestamp 1644511149
transform 1 0 34960 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_380
timestamp 1644511149
transform 1 0 36064 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_392
timestamp 1644511149
transform 1 0 37168 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_404
timestamp 1644511149
transform 1 0 38272 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_15
timestamp 1644511149
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_27
timestamp 1644511149
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_39
timestamp 1644511149
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1644511149
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1644511149
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_125
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_137
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_149
timestamp 1644511149
transform 1 0 14812 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_164
timestamp 1644511149
transform 1 0 16192 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_169
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_179
timestamp 1644511149
transform 1 0 17572 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_192
timestamp 1644511149
transform 1 0 18768 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_204
timestamp 1644511149
transform 1 0 19872 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_212
timestamp 1644511149
transform 1 0 20608 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_220
timestamp 1644511149
transform 1 0 21344 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_225
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_239
timestamp 1644511149
transform 1 0 23092 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_246
timestamp 1644511149
transform 1 0 23736 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_255
timestamp 1644511149
transform 1 0 24564 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_264
timestamp 1644511149
transform 1 0 25392 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_276
timestamp 1644511149
transform 1 0 26496 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_287
timestamp 1644511149
transform 1 0 27508 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_55_306
timestamp 1644511149
transform 1 0 29256 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_322
timestamp 1644511149
transform 1 0 30728 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_332
timestamp 1644511149
transform 1 0 31648 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_344
timestamp 1644511149
transform 1 0 32752 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_55_359
timestamp 1644511149
transform 1 0 34132 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_371
timestamp 1644511149
transform 1 0 35236 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_383
timestamp 1644511149
transform 1 0 36340 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1644511149
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_393
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_405
timestamp 1644511149
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_7
timestamp 1644511149
transform 1 0 1748 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_19
timestamp 1644511149
transform 1 0 2852 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1644511149
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_121
timestamp 1644511149
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1644511149
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1644511149
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_153
timestamp 1644511149
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_165
timestamp 1644511149
transform 1 0 16284 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_169
timestamp 1644511149
transform 1 0 16652 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_180
timestamp 1644511149
transform 1 0 17664 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_187
timestamp 1644511149
transform 1 0 18308 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1644511149
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_197
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_215
timestamp 1644511149
transform 1 0 20884 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_226
timestamp 1644511149
transform 1 0 21896 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_233
timestamp 1644511149
transform 1 0 22540 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_241
timestamp 1644511149
transform 1 0 23276 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_248
timestamp 1644511149
transform 1 0 23920 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_258
timestamp 1644511149
transform 1 0 24840 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_265
timestamp 1644511149
transform 1 0 25484 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_277
timestamp 1644511149
transform 1 0 26588 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_287
timestamp 1644511149
transform 1 0 27508 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_293
timestamp 1644511149
transform 1 0 28060 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_300
timestamp 1644511149
transform 1 0 28704 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_317
timestamp 1644511149
transform 1 0 30268 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_321
timestamp 1644511149
transform 1 0 30636 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_328
timestamp 1644511149
transform 1 0 31280 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_335
timestamp 1644511149
transform 1 0 31924 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_348
timestamp 1644511149
transform 1 0 33120 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_359
timestamp 1644511149
transform 1 0 34132 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1644511149
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_372
timestamp 1644511149
transform 1 0 35328 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_384
timestamp 1644511149
transform 1 0 36432 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_396
timestamp 1644511149
transform 1 0 37536 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_404
timestamp 1644511149
transform 1 0 38272 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1644511149
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_27
timestamp 1644511149
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_39
timestamp 1644511149
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1644511149
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1644511149
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_125
timestamp 1644511149
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_137
timestamp 1644511149
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_149
timestamp 1644511149
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1644511149
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1644511149
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_181
timestamp 1644511149
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_193
timestamp 1644511149
transform 1 0 18860 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_202
timestamp 1644511149
transform 1 0 19688 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_214
timestamp 1644511149
transform 1 0 20792 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_222
timestamp 1644511149
transform 1 0 21528 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_234
timestamp 1644511149
transform 1 0 22632 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_254
timestamp 1644511149
transform 1 0 24472 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_261
timestamp 1644511149
transform 1 0 25116 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_265
timestamp 1644511149
transform 1 0 25484 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_276
timestamp 1644511149
transform 1 0 26496 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_287
timestamp 1644511149
transform 1 0 27508 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_291
timestamp 1644511149
transform 1 0 27876 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_309
timestamp 1644511149
transform 1 0 29532 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_318
timestamp 1644511149
transform 1 0 30360 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_332
timestamp 1644511149
transform 1 0 31648 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_337
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_351
timestamp 1644511149
transform 1 0 33396 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_362
timestamp 1644511149
transform 1 0 34408 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_374
timestamp 1644511149
transform 1 0 35512 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_386
timestamp 1644511149
transform 1 0 36616 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_57_393
timestamp 1644511149
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_405
timestamp 1644511149
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1644511149
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1644511149
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_121
timestamp 1644511149
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1644511149
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_153
timestamp 1644511149
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_165
timestamp 1644511149
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_177
timestamp 1644511149
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1644511149
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1644511149
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_197
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_206
timestamp 1644511149
transform 1 0 20056 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_215
timestamp 1644511149
transform 1 0 20884 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_224
timestamp 1644511149
transform 1 0 21712 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_236
timestamp 1644511149
transform 1 0 22816 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_242
timestamp 1644511149
transform 1 0 23368 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_248
timestamp 1644511149
transform 1 0 23920 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_274
timestamp 1644511149
transform 1 0 26312 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_288
timestamp 1644511149
transform 1 0 27600 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_58_300
timestamp 1644511149
transform 1 0 28704 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_315
timestamp 1644511149
transform 1 0 30084 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_322
timestamp 1644511149
transform 1 0 30728 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_331
timestamp 1644511149
transform 1 0 31556 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_340
timestamp 1644511149
transform 1 0 32384 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_348
timestamp 1644511149
transform 1 0 33120 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_360
timestamp 1644511149
transform 1 0 34224 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_365
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_377
timestamp 1644511149
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_389
timestamp 1644511149
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_401
timestamp 1644511149
transform 1 0 37996 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1644511149
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1644511149
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1644511149
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1644511149
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1644511149
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_125
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_137
timestamp 1644511149
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_149
timestamp 1644511149
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1644511149
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1644511149
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_181
timestamp 1644511149
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_193
timestamp 1644511149
transform 1 0 18860 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_202
timestamp 1644511149
transform 1 0 19688 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_213
timestamp 1644511149
transform 1 0 20700 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_220
timestamp 1644511149
transform 1 0 21344 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_234
timestamp 1644511149
transform 1 0 22632 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_240
timestamp 1644511149
transform 1 0 23184 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_254
timestamp 1644511149
transform 1 0 24472 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_268
timestamp 1644511149
transform 1 0 25760 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_275
timestamp 1644511149
transform 1 0 26404 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1644511149
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_284
timestamp 1644511149
transform 1 0 27232 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_293
timestamp 1644511149
transform 1 0 28060 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_302
timestamp 1644511149
transform 1 0 28888 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_309
timestamp 1644511149
transform 1 0 29532 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_315
timestamp 1644511149
transform 1 0 30084 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_321
timestamp 1644511149
transform 1 0 30636 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_330
timestamp 1644511149
transform 1 0 31464 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_341
timestamp 1644511149
transform 1 0 32476 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_353
timestamp 1644511149
transform 1 0 33580 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_365
timestamp 1644511149
transform 1 0 34684 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_377
timestamp 1644511149
transform 1 0 35788 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_389
timestamp 1644511149
transform 1 0 36892 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_59_393
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_403
timestamp 1644511149
transform 1 0 38180 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1644511149
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1644511149
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1644511149
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1644511149
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_121
timestamp 1644511149
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_153
timestamp 1644511149
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_165
timestamp 1644511149
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_177
timestamp 1644511149
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1644511149
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1644511149
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_197
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_205
timestamp 1644511149
transform 1 0 19964 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_210
timestamp 1644511149
transform 1 0 20424 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_217
timestamp 1644511149
transform 1 0 21068 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_229
timestamp 1644511149
transform 1 0 22172 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_241
timestamp 1644511149
transform 1 0 23276 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_248
timestamp 1644511149
transform 1 0 23920 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_260
timestamp 1644511149
transform 1 0 25024 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_278
timestamp 1644511149
transform 1 0 26680 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_286
timestamp 1644511149
transform 1 0 27416 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_294
timestamp 1644511149
transform 1 0 28152 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1644511149
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1644511149
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_60_309
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_314
timestamp 1644511149
transform 1 0 29992 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_327
timestamp 1644511149
transform 1 0 31188 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_336
timestamp 1644511149
transform 1 0 32016 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_348
timestamp 1644511149
transform 1 0 33120 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_360
timestamp 1644511149
transform 1 0 34224 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_365
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_377
timestamp 1644511149
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_389
timestamp 1644511149
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_401
timestamp 1644511149
transform 1 0 37996 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1644511149
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_27
timestamp 1644511149
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_39
timestamp 1644511149
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1644511149
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1644511149
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_93
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1644511149
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_149
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1644511149
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1644511149
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_181
timestamp 1644511149
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_193
timestamp 1644511149
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_205
timestamp 1644511149
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1644511149
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1644511149
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_225
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_237
timestamp 1644511149
transform 1 0 22908 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_243
timestamp 1644511149
transform 1 0 23460 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_247
timestamp 1644511149
transform 1 0 23828 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_255
timestamp 1644511149
transform 1 0 24564 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_61_264
timestamp 1644511149
transform 1 0 25392 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_276
timestamp 1644511149
transform 1 0 26496 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_290
timestamp 1644511149
transform 1 0 27784 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_294
timestamp 1644511149
transform 1 0 28152 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_302
timestamp 1644511149
transform 1 0 28888 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_311
timestamp 1644511149
transform 1 0 29716 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_332
timestamp 1644511149
transform 1 0 31648 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_342
timestamp 1644511149
transform 1 0 32568 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_349
timestamp 1644511149
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_361
timestamp 1644511149
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_373
timestamp 1644511149
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1644511149
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1644511149
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_393
timestamp 1644511149
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1644511149
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_15
timestamp 1644511149
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1644511149
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1644511149
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1644511149
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_109
timestamp 1644511149
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_121
timestamp 1644511149
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1644511149
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1644511149
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_153
timestamp 1644511149
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_165
timestamp 1644511149
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_177
timestamp 1644511149
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1644511149
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1644511149
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_197
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_209
timestamp 1644511149
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_221
timestamp 1644511149
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_233
timestamp 1644511149
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_248
timestamp 1644511149
transform 1 0 23920 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_253
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_262
timestamp 1644511149
transform 1 0 25208 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_270
timestamp 1644511149
transform 1 0 25944 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_278
timestamp 1644511149
transform 1 0 26680 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_290
timestamp 1644511149
transform 1 0 27784 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_294
timestamp 1644511149
transform 1 0 28152 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_304
timestamp 1644511149
transform 1 0 29072 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_309
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_315
timestamp 1644511149
transform 1 0 30084 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_325
timestamp 1644511149
transform 1 0 31004 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_335
timestamp 1644511149
transform 1 0 31924 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_343
timestamp 1644511149
transform 1 0 32660 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_355
timestamp 1644511149
transform 1 0 33764 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1644511149
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_377
timestamp 1644511149
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_389
timestamp 1644511149
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_401
timestamp 1644511149
transform 1 0 37996 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1644511149
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_27
timestamp 1644511149
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_39
timestamp 1644511149
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1644511149
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1644511149
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1644511149
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1644511149
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_137
timestamp 1644511149
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_149
timestamp 1644511149
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1644511149
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1644511149
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_181
timestamp 1644511149
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_193
timestamp 1644511149
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_205
timestamp 1644511149
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1644511149
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1644511149
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_225
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_237
timestamp 1644511149
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_249
timestamp 1644511149
transform 1 0 24012 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_255
timestamp 1644511149
transform 1 0 24564 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_268
timestamp 1644511149
transform 1 0 25760 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_275
timestamp 1644511149
transform 1 0 26404 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1644511149
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_63_281
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_63_291
timestamp 1644511149
transform 1 0 27876 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_63_303
timestamp 1644511149
transform 1 0 28980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_309
timestamp 1644511149
transform 1 0 29532 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_313
timestamp 1644511149
transform 1 0 29900 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_324
timestamp 1644511149
transform 1 0 30912 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_337
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_349
timestamp 1644511149
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_361
timestamp 1644511149
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_373
timestamp 1644511149
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1644511149
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1644511149
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_393
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_405
timestamp 1644511149
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1644511149
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1644511149
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_33
timestamp 1644511149
transform 1 0 4140 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_45
timestamp 1644511149
transform 1 0 5244 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_53
timestamp 1644511149
transform 1 0 5980 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_57
timestamp 1644511149
transform 1 0 6348 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_69
timestamp 1644511149
transform 1 0 7452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_81
timestamp 1644511149
transform 1 0 8556 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_97
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_109
timestamp 1644511149
transform 1 0 11132 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_113
timestamp 1644511149
transform 1 0 11500 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_125
timestamp 1644511149
transform 1 0 12604 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_137
timestamp 1644511149
transform 1 0 13708 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_145
timestamp 1644511149
transform 1 0 14444 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_157
timestamp 1644511149
transform 1 0 15548 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_165
timestamp 1644511149
transform 1 0 16284 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_169
timestamp 1644511149
transform 1 0 16652 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_181
timestamp 1644511149
transform 1 0 17756 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_193
timestamp 1644511149
transform 1 0 18860 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_197
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_209
timestamp 1644511149
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_221
timestamp 1644511149
transform 1 0 21436 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_225
timestamp 1644511149
transform 1 0 21804 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_237
timestamp 1644511149
transform 1 0 22908 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_243
timestamp 1644511149
transform 1 0 23460 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_248
timestamp 1644511149
transform 1 0 23920 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_253
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_259
timestamp 1644511149
transform 1 0 24932 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_265
timestamp 1644511149
transform 1 0 25484 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_275
timestamp 1644511149
transform 1 0 26404 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_279
timestamp 1644511149
transform 1 0 26772 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_286
timestamp 1644511149
transform 1 0 27416 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_294
timestamp 1644511149
transform 1 0 28152 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1644511149
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1644511149
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_309
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_320
timestamp 1644511149
transform 1 0 30544 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_332
timestamp 1644511149
transform 1 0 31648 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_337
timestamp 1644511149
transform 1 0 32108 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_349
timestamp 1644511149
transform 1 0 33212 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_361
timestamp 1644511149
transform 1 0 34316 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_369
timestamp 1644511149
transform 1 0 35052 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_381
timestamp 1644511149
transform 1 0 36156 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_389
timestamp 1644511149
transform 1 0 36892 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_393
timestamp 1644511149
transform 1 0 37260 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_405
timestamp 1644511149
transform 1 0 38364 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0875_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16192 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0876_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18308 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0877_
timestamp 1644511149
transform 1 0 16100 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _0878_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14904 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0879_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0880_
timestamp 1644511149
transform 1 0 17480 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0881_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15916 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0882_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18032 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0883_
timestamp 1644511149
transform 1 0 17848 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0884_
timestamp 1644511149
transform 1 0 18676 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0885_
timestamp 1644511149
transform 1 0 16192 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__and3b_1  _0886_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16284 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0887_
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0888_
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0889_
timestamp 1644511149
transform 1 0 23368 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0890_
timestamp 1644511149
transform 1 0 24656 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0891_
timestamp 1644511149
transform 1 0 26680 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0892_
timestamp 1644511149
transform 1 0 25944 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0893_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16192 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0894_
timestamp 1644511149
transform 1 0 22724 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0895_
timestamp 1644511149
transform 1 0 24748 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _0896_
timestamp 1644511149
transform 1 0 15456 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0897_
timestamp 1644511149
transform 1 0 18124 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_2  _0898_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22264 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0899_
timestamp 1644511149
transform 1 0 15916 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0900_
timestamp 1644511149
transform 1 0 20700 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0901_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22356 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_1  _0902_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21252 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  _0903_
timestamp 1644511149
transform 1 0 18860 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0904_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19228 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or3_2  _0905_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16744 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0906_
timestamp 1644511149
transform 1 0 17664 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _0907_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17664 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0908_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21068 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0909_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19688 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0910_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18308 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0911_
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _0912_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17756 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0913_
timestamp 1644511149
transform 1 0 20700 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0914_
timestamp 1644511149
transform 1 0 19964 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0915_
timestamp 1644511149
transform 1 0 20976 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0916_
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0917_
timestamp 1644511149
transform 1 0 21804 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0918_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16928 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0919_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16928 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0920_
timestamp 1644511149
transform 1 0 16100 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0921_
timestamp 1644511149
transform 1 0 21804 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0922_
timestamp 1644511149
transform 1 0 20976 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a311o_1  _0923_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20424 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0924_
timestamp 1644511149
transform 1 0 20700 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0925_
timestamp 1644511149
transform 1 0 18492 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _0926_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19688 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0927_
timestamp 1644511149
transform 1 0 20148 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0928_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19412 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0929_
timestamp 1644511149
transform 1 0 19780 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0930_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16928 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0931_
timestamp 1644511149
transform 1 0 16376 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _0932_
timestamp 1644511149
transform 1 0 15548 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0933_
timestamp 1644511149
transform 1 0 22908 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0934_
timestamp 1644511149
transform 1 0 22172 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_2  _0935_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19412 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _0936_
timestamp 1644511149
transform 1 0 19780 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0937_
timestamp 1644511149
transform 1 0 19964 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0938_
timestamp 1644511149
transform 1 0 18768 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0939_
timestamp 1644511149
transform 1 0 20976 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0940_
timestamp 1644511149
transform 1 0 18952 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0941_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15548 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_2  _0942_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16284 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0943_
timestamp 1644511149
transform 1 0 15732 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0944_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15180 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0945_
timestamp 1644511149
transform 1 0 15916 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0946_
timestamp 1644511149
transform 1 0 18308 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_2  _0947_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20792 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_2  _0948_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16744 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0949_
timestamp 1644511149
transform 1 0 15916 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0950_
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0951_
timestamp 1644511149
transform 1 0 15088 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0952_
timestamp 1644511149
transform 1 0 15272 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0953_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15548 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0954_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16744 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o31ai_2  _0955_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16744 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0956_
timestamp 1644511149
transform 1 0 17756 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _0957_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19136 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a311oi_4  _0958_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_2  _0959_
timestamp 1644511149
transform 1 0 17480 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o31ai_2  _0960_
timestamp 1644511149
transform 1 0 17664 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _0961_
timestamp 1644511149
transform 1 0 18308 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0962_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18216 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0963_
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0964_
timestamp 1644511149
transform 1 0 17940 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0965_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19596 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0966_
timestamp 1644511149
transform 1 0 21068 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0967_
timestamp 1644511149
transform 1 0 20332 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0968_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20056 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0969_
timestamp 1644511149
transform 1 0 21252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0970_
timestamp 1644511149
transform 1 0 20608 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0971_
timestamp 1644511149
transform 1 0 24104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0972_
timestamp 1644511149
transform 1 0 23828 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0973_
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0974_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19136 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_1  _0975_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20424 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0976_
timestamp 1644511149
transform 1 0 18032 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _0977_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16836 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _0978_
timestamp 1644511149
transform 1 0 23460 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0979_
timestamp 1644511149
transform 1 0 22264 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0980_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20332 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0981_
timestamp 1644511149
transform 1 0 21252 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _0982_
timestamp 1644511149
transform 1 0 20056 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0983_
timestamp 1644511149
transform 1 0 17940 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0984_
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0985_
timestamp 1644511149
transform 1 0 23460 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _0986_
timestamp 1644511149
transform 1 0 21712 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0987_
timestamp 1644511149
transform 1 0 17388 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0988_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23368 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0989_
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0990_
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0991_
timestamp 1644511149
transform 1 0 23460 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0992_
timestamp 1644511149
transform 1 0 23460 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0993_
timestamp 1644511149
transform 1 0 29992 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _0994_
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0995_
timestamp 1644511149
transform 1 0 21252 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0996_
timestamp 1644511149
transform 1 0 21068 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0997_
timestamp 1644511149
transform 1 0 20148 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0998_
timestamp 1644511149
transform 1 0 19412 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0999_
timestamp 1644511149
transform 1 0 20792 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1000_
timestamp 1644511149
transform 1 0 20056 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1001_
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1002_
timestamp 1644511149
transform 1 0 23644 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1003_
timestamp 1644511149
transform 1 0 28704 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1004_
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1005_
timestamp 1644511149
transform 1 0 24472 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1006_
timestamp 1644511149
transform 1 0 22816 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1007_
timestamp 1644511149
transform 1 0 22908 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_2  _1008_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23092 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_2  _1009_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28060 0 -1 32640
box -38 -48 1234 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1010_
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1011_
timestamp 1644511149
transform 1 0 31740 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1012_
timestamp 1644511149
transform 1 0 28244 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1013_
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1014_
timestamp 1644511149
transform 1 0 26036 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1015_
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1016_
timestamp 1644511149
transform 1 0 25668 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _1017_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26036 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1018_
timestamp 1644511149
transform 1 0 23460 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1019_
timestamp 1644511149
transform 1 0 23644 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1020_
timestamp 1644511149
transform 1 0 22172 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1021_
timestamp 1644511149
transform 1 0 24656 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1022_
timestamp 1644511149
transform 1 0 26128 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_4  _1023_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25116 0 -1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_1  _1024_
timestamp 1644511149
transform 1 0 27600 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1025_
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1026_
timestamp 1644511149
transform 1 0 28244 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_4  _1027_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27968 0 -1 33728
box -38 -48 1602 592
use sky130_fd_sc_hd__and3_1  _1028_
timestamp 1644511149
transform 1 0 20884 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _1029_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22356 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1030_
timestamp 1644511149
transform 1 0 24840 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a311oi_4  _1031_
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1032_
timestamp 1644511149
transform 1 0 26680 0 1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1033_
timestamp 1644511149
transform 1 0 23184 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1034_
timestamp 1644511149
transform 1 0 24932 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1035_
timestamp 1644511149
transform 1 0 24288 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1036_
timestamp 1644511149
transform 1 0 25208 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1037_
timestamp 1644511149
transform 1 0 25576 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _1038_
timestamp 1644511149
transform 1 0 27048 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1039_
timestamp 1644511149
transform 1 0 24840 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__o21a_1  _1040_
timestamp 1644511149
transform 1 0 28152 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1041_
timestamp 1644511149
transform 1 0 28428 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1042_
timestamp 1644511149
transform 1 0 27784 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1043_
timestamp 1644511149
transform 1 0 28152 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1044_
timestamp 1644511149
transform 1 0 28520 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1045_
timestamp 1644511149
transform 1 0 27508 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1046_
timestamp 1644511149
transform 1 0 27968 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1047_
timestamp 1644511149
transform 1 0 29256 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _1048_
timestamp 1644511149
transform 1 0 28244 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1049_
timestamp 1644511149
transform 1 0 30268 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _1050_
timestamp 1644511149
transform 1 0 23736 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1051_
timestamp 1644511149
transform 1 0 24932 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1052_
timestamp 1644511149
transform 1 0 26956 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1053_
timestamp 1644511149
transform 1 0 29256 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1054_
timestamp 1644511149
transform 1 0 29900 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1055_
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1056_
timestamp 1644511149
transform 1 0 29624 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1057_
timestamp 1644511149
transform 1 0 24288 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1058_
timestamp 1644511149
transform 1 0 29072 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1059_
timestamp 1644511149
transform 1 0 24932 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1060_
timestamp 1644511149
transform 1 0 25116 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1061_
timestamp 1644511149
transform 1 0 26128 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _1062_
timestamp 1644511149
transform 1 0 25484 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1063_
timestamp 1644511149
transform 1 0 31924 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1064_
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1065_
timestamp 1644511149
transform 1 0 29900 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1066_
timestamp 1644511149
transform 1 0 28152 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1067_
timestamp 1644511149
transform 1 0 33580 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1068_
timestamp 1644511149
transform 1 0 30452 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _1069_
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1070_
timestamp 1644511149
transform 1 0 33120 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1071_
timestamp 1644511149
transform 1 0 31832 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1072_
timestamp 1644511149
transform 1 0 30728 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1073_
timestamp 1644511149
transform 1 0 31096 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1074_
timestamp 1644511149
transform 1 0 30636 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1075_
timestamp 1644511149
transform 1 0 32936 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1076_
timestamp 1644511149
transform 1 0 33672 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1077_
timestamp 1644511149
transform 1 0 33396 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1078_
timestamp 1644511149
transform 1 0 33488 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1079_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32292 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1080_
timestamp 1644511149
transform 1 0 30176 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1081_
timestamp 1644511149
transform 1 0 31556 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1082_
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _1083_
timestamp 1644511149
transform 1 0 30452 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1084_
timestamp 1644511149
transform 1 0 30268 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1085_
timestamp 1644511149
transform 1 0 23552 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _1086_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23276 0 -1 34816
box -38 -48 1234 592
use sky130_fd_sc_hd__o21a_1  _1087_
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_2  _1088_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25760 0 1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _1089_
timestamp 1644511149
transform 1 0 25944 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _1090_
timestamp 1644511149
transform 1 0 25852 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1091_
timestamp 1644511149
transform 1 0 33580 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1092_
timestamp 1644511149
transform 1 0 24932 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1093_
timestamp 1644511149
transform 1 0 23644 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1094_
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1095_
timestamp 1644511149
transform 1 0 24748 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1096_
timestamp 1644511149
transform 1 0 24748 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1097_
timestamp 1644511149
transform 1 0 24196 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1098_
timestamp 1644511149
transform 1 0 26128 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1099_
timestamp 1644511149
transform 1 0 29624 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1100_
timestamp 1644511149
transform 1 0 29624 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1101_
timestamp 1644511149
transform 1 0 31372 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__o21bai_1  _1102_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25852 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _1103_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30820 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_2  _1104_
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1105_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30728 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1106_
timestamp 1644511149
transform 1 0 28244 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1107_
timestamp 1644511149
transform 1 0 31004 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1108_
timestamp 1644511149
transform 1 0 32292 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1109_
timestamp 1644511149
transform 1 0 32936 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1110_
timestamp 1644511149
transform 1 0 30360 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _1111_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28060 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1112_
timestamp 1644511149
transform 1 0 28704 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1113_
timestamp 1644511149
transform 1 0 32476 0 -1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _1114_
timestamp 1644511149
transform 1 0 31648 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1115_
timestamp 1644511149
transform 1 0 32752 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1116_
timestamp 1644511149
transform 1 0 31096 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1117_
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1118_
timestamp 1644511149
transform 1 0 24748 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1119_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30912 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1120_
timestamp 1644511149
transform 1 0 31096 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1121_
timestamp 1644511149
transform 1 0 30268 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1122_
timestamp 1644511149
transform 1 0 33764 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1123_
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1124_
timestamp 1644511149
transform 1 0 33304 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _1125_
timestamp 1644511149
transform 1 0 30912 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1126_
timestamp 1644511149
transform 1 0 32292 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1127_
timestamp 1644511149
transform 1 0 30360 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1128_
timestamp 1644511149
transform 1 0 31372 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1129_
timestamp 1644511149
transform 1 0 33304 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1130_
timestamp 1644511149
transform 1 0 35144 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1131_
timestamp 1644511149
transform 1 0 28704 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1132_
timestamp 1644511149
transform 1 0 29532 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1133_
timestamp 1644511149
transform 1 0 31280 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1134_
timestamp 1644511149
transform 1 0 32568 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1135_
timestamp 1644511149
transform 1 0 32016 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1136_
timestamp 1644511149
transform 1 0 30544 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1137_
timestamp 1644511149
transform 1 0 29716 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _1138_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 31096 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _1139_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29992 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1140_
timestamp 1644511149
transform 1 0 25760 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1141_
timestamp 1644511149
transform 1 0 25944 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1142_
timestamp 1644511149
transform 1 0 26956 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1143_
timestamp 1644511149
transform 1 0 28428 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1144_
timestamp 1644511149
transform 1 0 27232 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1145_
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1146_
timestamp 1644511149
transform 1 0 26128 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _1147_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28244 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__o22ai_1  _1148_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25024 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1149_
timestamp 1644511149
transform 1 0 24932 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1150_
timestamp 1644511149
transform 1 0 23920 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o22ai_2  _1151_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25576 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1152_
timestamp 1644511149
transform 1 0 25576 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1153_
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1154_
timestamp 1644511149
transform 1 0 26680 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1155_
timestamp 1644511149
transform 1 0 25392 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1156_
timestamp 1644511149
transform 1 0 26128 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1157_
timestamp 1644511149
transform 1 0 26036 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1158_
timestamp 1644511149
transform 1 0 32476 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1159_
timestamp 1644511149
transform 1 0 32292 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1160_
timestamp 1644511149
transform 1 0 25668 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1161_
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1162_
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1163_
timestamp 1644511149
transform 1 0 26864 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1164_
timestamp 1644511149
transform 1 0 13248 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1165_
timestamp 1644511149
transform 1 0 20884 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1166_
timestamp 1644511149
transform 1 0 25852 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1167_
timestamp 1644511149
transform 1 0 15824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1168_
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1169_
timestamp 1644511149
transform 1 0 17940 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1170_
timestamp 1644511149
transform 1 0 24748 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1171_
timestamp 1644511149
transform 1 0 23460 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1172_
timestamp 1644511149
transform 1 0 24104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1173_
timestamp 1644511149
transform 1 0 24748 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1174_
timestamp 1644511149
transform 1 0 29624 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1175_
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1176_
timestamp 1644511149
transform 1 0 29164 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1177_
timestamp 1644511149
transform 1 0 28336 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1178_
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1179_
timestamp 1644511149
transform 1 0 26772 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1180_
timestamp 1644511149
transform 1 0 31188 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1181_
timestamp 1644511149
transform 1 0 31188 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1182_
timestamp 1644511149
transform 1 0 29624 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1183_
timestamp 1644511149
transform 1 0 28796 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1184_
timestamp 1644511149
transform 1 0 30176 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1185_
timestamp 1644511149
transform 1 0 27876 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1186_
timestamp 1644511149
transform 1 0 24748 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1187_
timestamp 1644511149
transform 1 0 28520 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1188_
timestamp 1644511149
transform 1 0 27416 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1189_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26864 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1190_
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1191_
timestamp 1644511149
transform 1 0 24196 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1192_
timestamp 1644511149
transform 1 0 24840 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1193_
timestamp 1644511149
transform 1 0 24012 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1194_
timestamp 1644511149
transform 1 0 24564 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1195_
timestamp 1644511149
transform 1 0 29992 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1196_
timestamp 1644511149
transform 1 0 31096 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1197_
timestamp 1644511149
transform 1 0 30268 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1198_
timestamp 1644511149
transform 1 0 30544 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1199_
timestamp 1644511149
transform 1 0 30636 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1200_
timestamp 1644511149
transform 1 0 30636 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1201_
timestamp 1644511149
transform 1 0 30544 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1202_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30544 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1203_
timestamp 1644511149
transform 1 0 30636 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1204_
timestamp 1644511149
transform 1 0 30820 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1205_
timestamp 1644511149
transform 1 0 30452 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1206_
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1207_
timestamp 1644511149
transform 1 0 28704 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1208_
timestamp 1644511149
transform 1 0 29808 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1209_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28336 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1210_
timestamp 1644511149
transform 1 0 26128 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _1211_
timestamp 1644511149
transform 1 0 29348 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1212_
timestamp 1644511149
transform 1 0 28060 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1213_
timestamp 1644511149
transform 1 0 28060 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1214_
timestamp 1644511149
transform 1 0 27508 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1215_
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1216_
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1217_
timestamp 1644511149
transform 1 0 21804 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__o311a_1  _1218_
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _1219_
timestamp 1644511149
transform 1 0 29900 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_4  _1220_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27968 0 -1 25024
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_2  _1221_
timestamp 1644511149
transform 1 0 28980 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _1222_
timestamp 1644511149
transform 1 0 28060 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1223_
timestamp 1644511149
transform 1 0 27692 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1224_
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1225_
timestamp 1644511149
transform 1 0 32752 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1226_
timestamp 1644511149
transform 1 0 30176 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _1227_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30636 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1228_
timestamp 1644511149
transform 1 0 30912 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1229_
timestamp 1644511149
transform 1 0 30268 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1230_
timestamp 1644511149
transform 1 0 30544 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1231_
timestamp 1644511149
transform 1 0 31556 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1232_
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1233_
timestamp 1644511149
transform 1 0 32384 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1234_
timestamp 1644511149
transform 1 0 31188 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1235_
timestamp 1644511149
transform 1 0 31464 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1236_
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1237_
timestamp 1644511149
transform 1 0 31280 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1238_
timestamp 1644511149
transform 1 0 30636 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1239_
timestamp 1644511149
transform 1 0 29440 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1240_
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1241_
timestamp 1644511149
transform 1 0 27048 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1242_
timestamp 1644511149
transform 1 0 22356 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_1  _1243_
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1244_
timestamp 1644511149
transform 1 0 22632 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1245_
timestamp 1644511149
transform 1 0 31740 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1246_
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1247_
timestamp 1644511149
transform 1 0 22448 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1248_
timestamp 1644511149
transform 1 0 26404 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1249_
timestamp 1644511149
transform 1 0 32384 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1250_
timestamp 1644511149
transform 1 0 32292 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1251_
timestamp 1644511149
transform 1 0 32200 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1252_
timestamp 1644511149
transform 1 0 32660 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1253_
timestamp 1644511149
transform 1 0 29348 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1254_
timestamp 1644511149
transform 1 0 29808 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1255_
timestamp 1644511149
transform 1 0 30268 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1256_
timestamp 1644511149
transform 1 0 31188 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1257_
timestamp 1644511149
transform 1 0 31464 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1258_
timestamp 1644511149
transform 1 0 33028 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1259_
timestamp 1644511149
transform 1 0 32752 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1260_
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1261_
timestamp 1644511149
transform 1 0 32752 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_2  _1262_
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1263_
timestamp 1644511149
transform 1 0 33212 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand3b_1  _1264_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32936 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1265_
timestamp 1644511149
transform 1 0 32660 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1266_
timestamp 1644511149
transform 1 0 33764 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1267_
timestamp 1644511149
transform 1 0 32936 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1268_
timestamp 1644511149
transform 1 0 32200 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1269_
timestamp 1644511149
transform 1 0 27508 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1270_
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1271_
timestamp 1644511149
transform 1 0 26864 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1272_
timestamp 1644511149
transform 1 0 27600 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1273_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28520 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1274_
timestamp 1644511149
transform 1 0 28336 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _1275_
timestamp 1644511149
transform 1 0 27968 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1276_
timestamp 1644511149
transform 1 0 27876 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1277_
timestamp 1644511149
transform 1 0 28244 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1278_
timestamp 1644511149
transform 1 0 27232 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1279_
timestamp 1644511149
transform 1 0 27140 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1280_
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_1  _1281_
timestamp 1644511149
transform 1 0 28704 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _1282_
timestamp 1644511149
transform 1 0 25760 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _1283_
timestamp 1644511149
transform 1 0 26128 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1284_
timestamp 1644511149
transform 1 0 26588 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1285_
timestamp 1644511149
transform 1 0 25484 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _1286_
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1287_
timestamp 1644511149
transform 1 0 23000 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1288_
timestamp 1644511149
transform 1 0 24012 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1289_
timestamp 1644511149
transform 1 0 25760 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1290_
timestamp 1644511149
transform 1 0 24472 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1291_
timestamp 1644511149
transform 1 0 25116 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1292_
timestamp 1644511149
transform 1 0 26588 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1293_
timestamp 1644511149
transform 1 0 25484 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1294_
timestamp 1644511149
transform 1 0 26036 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1295_
timestamp 1644511149
transform 1 0 33580 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1296_
timestamp 1644511149
transform 1 0 27324 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _1297_
timestamp 1644511149
transform 1 0 33304 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1298_
timestamp 1644511149
transform 1 0 32476 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _1299_
timestamp 1644511149
transform 1 0 33672 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  _1300_
timestamp 1644511149
transform 1 0 34316 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _1301_
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1302_
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_2  _1303_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30360 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1304_
timestamp 1644511149
transform 1 0 33304 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1305_
timestamp 1644511149
transform 1 0 29440 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1306_
timestamp 1644511149
transform 1 0 29808 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1307_
timestamp 1644511149
transform 1 0 33672 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1308_
timestamp 1644511149
transform 1 0 34316 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1309_
timestamp 1644511149
transform 1 0 35328 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1310_
timestamp 1644511149
transform 1 0 34868 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1311_
timestamp 1644511149
transform 1 0 35420 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1312_
timestamp 1644511149
transform 1 0 34408 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1313_
timestamp 1644511149
transform 1 0 33580 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1314_
timestamp 1644511149
transform 1 0 33672 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _1315_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1316_
timestamp 1644511149
transform 1 0 33120 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1317_
timestamp 1644511149
transform 1 0 34500 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1318_
timestamp 1644511149
transform 1 0 34776 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1319_
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1320_
timestamp 1644511149
transform 1 0 33764 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1321_
timestamp 1644511149
transform 1 0 25576 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1322_
timestamp 1644511149
transform 1 0 26864 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1323_
timestamp 1644511149
transform 1 0 25668 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1324_
timestamp 1644511149
transform 1 0 23552 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o311a_1  _1325_
timestamp 1644511149
transform 1 0 23736 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1326_
timestamp 1644511149
transform 1 0 24196 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1327_
timestamp 1644511149
transform 1 0 28244 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1328_
timestamp 1644511149
transform 1 0 22540 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1329_
timestamp 1644511149
transform 1 0 24196 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1330_
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__a21oi_1  _1331_
timestamp 1644511149
transform 1 0 25668 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1332_
timestamp 1644511149
transform 1 0 23000 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1333_
timestamp 1644511149
transform 1 0 33856 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1334_
timestamp 1644511149
transform 1 0 34776 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1335_
timestamp 1644511149
transform 1 0 35788 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1336_
timestamp 1644511149
transform 1 0 35880 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1337_
timestamp 1644511149
transform 1 0 35880 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _1338_
timestamp 1644511149
transform 1 0 35328 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1339_
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1340_
timestamp 1644511149
transform 1 0 28244 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _1341_
timestamp 1644511149
transform 1 0 33120 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_2  _1342_
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _1343_
timestamp 1644511149
transform 1 0 33488 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1344_
timestamp 1644511149
transform 1 0 35420 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1345_
timestamp 1644511149
transform 1 0 32844 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1346_
timestamp 1644511149
transform 1 0 33948 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1347_
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1348_
timestamp 1644511149
transform 1 0 22356 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1349_
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1350_
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1351_
timestamp 1644511149
transform 1 0 31924 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1352_
timestamp 1644511149
transform 1 0 35328 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1353_
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1354_
timestamp 1644511149
transform 1 0 34684 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1355_
timestamp 1644511149
transform 1 0 35512 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1356_
timestamp 1644511149
transform 1 0 35880 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1357_
timestamp 1644511149
transform 1 0 35788 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1358_
timestamp 1644511149
transform 1 0 36524 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1359_
timestamp 1644511149
transform 1 0 36248 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1360_
timestamp 1644511149
transform 1 0 35696 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1361_
timestamp 1644511149
transform 1 0 36064 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1362_
timestamp 1644511149
transform 1 0 35328 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o211ai_2  _1363_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 35604 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__a211o_1  _1364_
timestamp 1644511149
transform 1 0 35420 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _1365_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 34868 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__o2bb2a_1  _1366_
timestamp 1644511149
transform 1 0 34868 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1367_
timestamp 1644511149
transform 1 0 36156 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1368_
timestamp 1644511149
transform 1 0 34224 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1369_
timestamp 1644511149
transform 1 0 33120 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1370_
timestamp 1644511149
transform 1 0 25392 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1371_
timestamp 1644511149
transform 1 0 23184 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_2  _1372_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_1  _1373_
timestamp 1644511149
transform 1 0 32384 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _1374_
timestamp 1644511149
transform 1 0 23368 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1375_
timestamp 1644511149
transform 1 0 23092 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_2  _1376_
timestamp 1644511149
transform 1 0 22724 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _1377_
timestamp 1644511149
transform 1 0 21896 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1378_
timestamp 1644511149
transform 1 0 23368 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1379_
timestamp 1644511149
transform 1 0 23276 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1380_
timestamp 1644511149
transform 1 0 23552 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _1381_
timestamp 1644511149
transform 1 0 36616 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1382_
timestamp 1644511149
transform 1 0 37076 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1383_
timestamp 1644511149
transform 1 0 34316 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1384_
timestamp 1644511149
transform 1 0 34684 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1385_
timestamp 1644511149
transform 1 0 35696 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1386_
timestamp 1644511149
transform 1 0 36064 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1387_
timestamp 1644511149
transform 1 0 34316 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1388_
timestamp 1644511149
transform 1 0 28520 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1389_
timestamp 1644511149
transform 1 0 27140 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1390_
timestamp 1644511149
transform 1 0 27416 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_2  _1391_
timestamp 1644511149
transform 1 0 27508 0 1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _1392_
timestamp 1644511149
transform 1 0 34960 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1393_
timestamp 1644511149
transform 1 0 36432 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1394_
timestamp 1644511149
transform 1 0 30820 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1395_
timestamp 1644511149
transform 1 0 32936 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1396_
timestamp 1644511149
transform 1 0 33120 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1397_
timestamp 1644511149
transform 1 0 33948 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _1398_
timestamp 1644511149
transform 1 0 34868 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1399_
timestamp 1644511149
transform 1 0 35052 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1400_
timestamp 1644511149
transform 1 0 36064 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1401_
timestamp 1644511149
transform 1 0 36800 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1402_
timestamp 1644511149
transform 1 0 36432 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1403_
timestamp 1644511149
transform 1 0 37720 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1404_
timestamp 1644511149
transform 1 0 37444 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1405_
timestamp 1644511149
transform 1 0 37720 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1406_
timestamp 1644511149
transform 1 0 37168 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1407_
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1408_
timestamp 1644511149
transform 1 0 36432 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1409_
timestamp 1644511149
transform 1 0 34868 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1410_
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1411_
timestamp 1644511149
transform 1 0 21068 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1412_
timestamp 1644511149
transform 1 0 23552 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1413_
timestamp 1644511149
transform 1 0 23276 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_1  _1414_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22080 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1415_
timestamp 1644511149
transform 1 0 24288 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1416_
timestamp 1644511149
transform 1 0 30544 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1417_
timestamp 1644511149
transform 1 0 23092 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1418_
timestamp 1644511149
transform 1 0 35420 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1419_
timestamp 1644511149
transform 1 0 27416 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1420_
timestamp 1644511149
transform 1 0 33948 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1421_
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1422_
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1423_
timestamp 1644511149
transform 1 0 34316 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1424_
timestamp 1644511149
transform 1 0 35328 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1425_
timestamp 1644511149
transform 1 0 35696 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1426_
timestamp 1644511149
transform 1 0 28152 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1427_
timestamp 1644511149
transform 1 0 27416 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1428_
timestamp 1644511149
transform 1 0 26496 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1429_
timestamp 1644511149
transform 1 0 27232 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _1430_
timestamp 1644511149
transform 1 0 27140 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1431_
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1432_
timestamp 1644511149
transform 1 0 36984 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_1  _1433_
timestamp 1644511149
transform 1 0 37444 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _1434_
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1435_
timestamp 1644511149
transform 1 0 36064 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1436_
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1437_
timestamp 1644511149
transform 1 0 37536 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1438_
timestamp 1644511149
transform 1 0 36340 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1439_
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a221oi_1  _1440_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1441_
timestamp 1644511149
transform 1 0 31924 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1442_
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1443_
timestamp 1644511149
transform 1 0 37260 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1444_
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1445_
timestamp 1644511149
transform 1 0 36984 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _1446_
timestamp 1644511149
transform 1 0 21068 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1447_
timestamp 1644511149
transform 1 0 20332 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1448_
timestamp 1644511149
transform 1 0 20424 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _1449_
timestamp 1644511149
transform 1 0 25668 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1450_
timestamp 1644511149
transform 1 0 26128 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1451_
timestamp 1644511149
transform 1 0 24656 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _1452_
timestamp 1644511149
transform 1 0 25208 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1453_
timestamp 1644511149
transform 1 0 25760 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1454_
timestamp 1644511149
transform 1 0 22632 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _1455_
timestamp 1644511149
transform 1 0 21988 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1456_
timestamp 1644511149
transform 1 0 21436 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1457_
timestamp 1644511149
transform 1 0 20792 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1458_
timestamp 1644511149
transform 1 0 13984 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1459_
timestamp 1644511149
transform 1 0 19044 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1460_
timestamp 1644511149
transform 1 0 14720 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1461_
timestamp 1644511149
transform 1 0 20056 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1462_
timestamp 1644511149
transform 1 0 13248 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1463_
timestamp 1644511149
transform 1 0 18860 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1464_
timestamp 1644511149
transform 1 0 15456 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1465_
timestamp 1644511149
transform 1 0 14812 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor3b_1  _1466_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1467_
timestamp 1644511149
transform 1 0 17572 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1468_
timestamp 1644511149
transform 1 0 16560 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1469_
timestamp 1644511149
transform 1 0 13800 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1470_
timestamp 1644511149
transform 1 0 19872 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1471_
timestamp 1644511149
transform 1 0 11868 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1472_
timestamp 1644511149
transform 1 0 17848 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1473_
timestamp 1644511149
transform 1 0 10396 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1474_
timestamp 1644511149
transform 1 0 19964 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1475_
timestamp 1644511149
transform 1 0 8280 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1476_
timestamp 1644511149
transform 1 0 22448 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1477_
timestamp 1644511149
transform 1 0 23000 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1478_
timestamp 1644511149
transform 1 0 25392 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _1479_
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1480_
timestamp 1644511149
transform 1 0 28060 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1481_
timestamp 1644511149
transform 1 0 23552 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _1482_
timestamp 1644511149
transform 1 0 24932 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1483_
timestamp 1644511149
transform 1 0 24472 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1484_
timestamp 1644511149
transform 1 0 27232 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1485_
timestamp 1644511149
transform 1 0 25300 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1486_
timestamp 1644511149
transform 1 0 27324 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1487_
timestamp 1644511149
transform 1 0 25852 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1488_
timestamp 1644511149
transform 1 0 21712 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1489_
timestamp 1644511149
transform 1 0 23644 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _1490_
timestamp 1644511149
transform 1 0 22908 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1491_
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1492_
timestamp 1644511149
transform 1 0 24656 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1493_
timestamp 1644511149
transform 1 0 23552 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and2_2  _1494_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22724 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1495_
timestamp 1644511149
transform 1 0 23460 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1496_
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_2  _1497_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _1498_
timestamp 1644511149
transform 1 0 24840 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1499_
timestamp 1644511149
transform 1 0 27048 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1500_
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1501_
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _1502_
timestamp 1644511149
transform 1 0 28152 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1503_
timestamp 1644511149
transform 1 0 24288 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1504_
timestamp 1644511149
transform 1 0 24932 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1505_
timestamp 1644511149
transform 1 0 25852 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_2  _1506_
timestamp 1644511149
transform 1 0 25760 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1507_
timestamp 1644511149
transform 1 0 27600 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o221ai_4  _1508_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25484 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  _1509_
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _1510_
timestamp 1644511149
transform 1 0 23736 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _1511_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23368 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1512_
timestamp 1644511149
transform 1 0 25852 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _1513_
timestamp 1644511149
transform 1 0 25760 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_4  _1514_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25576 0 1 13056
box -38 -48 1326 592
use sky130_fd_sc_hd__a211o_1  _1515_
timestamp 1644511149
transform 1 0 26036 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1516_
timestamp 1644511149
transform 1 0 18216 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1517_
timestamp 1644511149
transform 1 0 15548 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1518_
timestamp 1644511149
transform 1 0 15916 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1519_
timestamp 1644511149
transform 1 0 15732 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1520_
timestamp 1644511149
transform 1 0 15732 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1521_
timestamp 1644511149
transform 1 0 14904 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1522_
timestamp 1644511149
transform 1 0 15088 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1523_
timestamp 1644511149
transform 1 0 14260 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1524_
timestamp 1644511149
transform 1 0 14168 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1525_
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1526_
timestamp 1644511149
transform 1 0 13340 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1527_
timestamp 1644511149
transform 1 0 14444 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1528_
timestamp 1644511149
transform 1 0 14996 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1529_
timestamp 1644511149
transform 1 0 13800 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1530_
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1531_
timestamp 1644511149
transform 1 0 13156 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1532_
timestamp 1644511149
transform 1 0 16560 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1533_
timestamp 1644511149
transform 1 0 13340 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1534_
timestamp 1644511149
transform 1 0 19044 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1535_
timestamp 1644511149
transform 1 0 20056 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1536_
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1537_
timestamp 1644511149
transform 1 0 20700 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1538_
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1539_
timestamp 1644511149
transform 1 0 18492 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1540_
timestamp 1644511149
transform 1 0 18308 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1541_
timestamp 1644511149
transform 1 0 19412 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1542_
timestamp 1644511149
transform 1 0 19780 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1543_
timestamp 1644511149
transform 1 0 17572 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1544_
timestamp 1644511149
transform 1 0 18400 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1545_
timestamp 1644511149
transform 1 0 18952 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1546_
timestamp 1644511149
transform 1 0 20056 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1547_
timestamp 1644511149
transform 1 0 17480 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1548_
timestamp 1644511149
transform 1 0 18492 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1549_
timestamp 1644511149
transform 1 0 19780 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1550_
timestamp 1644511149
transform 1 0 22908 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1551_
timestamp 1644511149
transform 1 0 20700 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1552_
timestamp 1644511149
transform 1 0 18860 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1553_
timestamp 1644511149
transform 1 0 19228 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1554_
timestamp 1644511149
transform 1 0 18492 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1555_
timestamp 1644511149
transform 1 0 18492 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1556_
timestamp 1644511149
transform 1 0 15272 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1557_
timestamp 1644511149
transform 1 0 17480 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1558_
timestamp 1644511149
transform 1 0 17756 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  _1559_
timestamp 1644511149
transform 1 0 15548 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1560_
timestamp 1644511149
transform 1 0 12788 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1561_
timestamp 1644511149
transform 1 0 12972 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1562_
timestamp 1644511149
transform 1 0 13340 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1563_
timestamp 1644511149
transform 1 0 12144 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1564_
timestamp 1644511149
transform 1 0 11500 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1565_
timestamp 1644511149
transform 1 0 11408 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1566_
timestamp 1644511149
transform 1 0 13064 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1567_
timestamp 1644511149
transform 1 0 13248 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1568_
timestamp 1644511149
transform 1 0 12512 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1569_
timestamp 1644511149
transform 1 0 14168 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1570_
timestamp 1644511149
transform 1 0 15916 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1571_
timestamp 1644511149
transform 1 0 13156 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1572_
timestamp 1644511149
transform 1 0 12512 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1573_
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1574_
timestamp 1644511149
transform 1 0 14076 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1575_
timestamp 1644511149
transform 1 0 13156 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1576_
timestamp 1644511149
transform 1 0 14904 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1577_
timestamp 1644511149
transform 1 0 15732 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1578_
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1579_
timestamp 1644511149
transform 1 0 15180 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1580_
timestamp 1644511149
transform 1 0 13800 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1581_
timestamp 1644511149
transform 1 0 13340 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1582_
timestamp 1644511149
transform 1 0 12052 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1583_
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1584_
timestamp 1644511149
transform 1 0 13340 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1585_
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1586_
timestamp 1644511149
transform 1 0 12328 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1587_
timestamp 1644511149
transform 1 0 9200 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1588_
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1589_
timestamp 1644511149
transform 1 0 14076 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1590_
timestamp 1644511149
transform 1 0 13156 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1591_
timestamp 1644511149
transform 1 0 12328 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1592_
timestamp 1644511149
transform 1 0 10856 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1593_
timestamp 1644511149
transform 1 0 11040 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1594_
timestamp 1644511149
transform 1 0 12788 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1595_
timestamp 1644511149
transform 1 0 11960 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1596_
timestamp 1644511149
transform 1 0 11868 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _1597_
timestamp 1644511149
transform 1 0 12788 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1598_
timestamp 1644511149
transform 1 0 10120 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1599_
timestamp 1644511149
transform 1 0 10120 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1600_
timestamp 1644511149
transform 1 0 12420 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1601_
timestamp 1644511149
transform 1 0 10028 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1602_
timestamp 1644511149
transform 1 0 11868 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1603_
timestamp 1644511149
transform 1 0 11408 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1604_
timestamp 1644511149
transform 1 0 12420 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1605_
timestamp 1644511149
transform 1 0 13432 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1606_
timestamp 1644511149
transform 1 0 11592 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1607_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11960 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1608_
timestamp 1644511149
transform 1 0 12144 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1609_
timestamp 1644511149
transform 1 0 12236 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1610_
timestamp 1644511149
transform 1 0 13248 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1611_
timestamp 1644511149
transform 1 0 12696 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1612_
timestamp 1644511149
transform 1 0 10580 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1613_
timestamp 1644511149
transform 1 0 9476 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1614_
timestamp 1644511149
transform 1 0 11132 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1615_
timestamp 1644511149
transform 1 0 14168 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1616_
timestamp 1644511149
transform 1 0 10120 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1617_
timestamp 1644511149
transform 1 0 11224 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1618_
timestamp 1644511149
transform 1 0 10488 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1619_
timestamp 1644511149
transform 1 0 10120 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1620_
timestamp 1644511149
transform 1 0 9384 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1621_
timestamp 1644511149
transform 1 0 9384 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1622_
timestamp 1644511149
transform 1 0 9936 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1623_
timestamp 1644511149
transform 1 0 10120 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1624_
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1625_
timestamp 1644511149
transform 1 0 9292 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1626_
timestamp 1644511149
transform 1 0 9568 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1627_
timestamp 1644511149
transform 1 0 9016 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1628_
timestamp 1644511149
transform 1 0 10488 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1629_
timestamp 1644511149
transform 1 0 9936 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1630_
timestamp 1644511149
transform 1 0 8556 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1631_
timestamp 1644511149
transform 1 0 8096 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_1  _1632_
timestamp 1644511149
transform 1 0 7728 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1633_
timestamp 1644511149
transform 1 0 8464 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1634_
timestamp 1644511149
transform 1 0 7544 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1635_
timestamp 1644511149
transform 1 0 8096 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1636_
timestamp 1644511149
transform 1 0 20884 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1637_
timestamp 1644511149
transform 1 0 19596 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1638_
timestamp 1644511149
transform 1 0 19136 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1639_
timestamp 1644511149
transform 1 0 21068 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1640_
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1641_
timestamp 1644511149
transform 1 0 19964 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1642_
timestamp 1644511149
transform 1 0 20792 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1643_
timestamp 1644511149
transform 1 0 18492 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1644_
timestamp 1644511149
transform 1 0 17848 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1645_
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1646_
timestamp 1644511149
transform 1 0 20332 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1647_
timestamp 1644511149
transform 1 0 20056 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1648_
timestamp 1644511149
transform 1 0 19688 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1649_
timestamp 1644511149
transform 1 0 17020 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _1650_
timestamp 1644511149
transform 1 0 17940 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1651_
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1652_
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1653_
timestamp 1644511149
transform 1 0 21988 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1654_
timestamp 1644511149
transform 1 0 21896 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1655_
timestamp 1644511149
transform 1 0 20792 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1656_
timestamp 1644511149
transform 1 0 22172 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1657_
timestamp 1644511149
transform 1 0 22724 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1658_
timestamp 1644511149
transform 1 0 21896 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1659_
timestamp 1644511149
transform 1 0 22356 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1660_
timestamp 1644511149
transform 1 0 23368 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1661_
timestamp 1644511149
transform 1 0 23184 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1662_
timestamp 1644511149
transform 1 0 12236 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1663_
timestamp 1644511149
transform 1 0 10764 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1664_
timestamp 1644511149
transform 1 0 16008 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1665_
timestamp 1644511149
transform 1 0 15732 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1666_
timestamp 1644511149
transform 1 0 14168 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1667_
timestamp 1644511149
transform 1 0 15088 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1668_
timestamp 1644511149
transform 1 0 17664 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1669_
timestamp 1644511149
transform 1 0 16192 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1670_
timestamp 1644511149
transform 1 0 17388 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1671_
timestamp 1644511149
transform 1 0 16836 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1672_
timestamp 1644511149
transform 1 0 16836 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1673_
timestamp 1644511149
transform 1 0 21068 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1674_
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1675_
timestamp 1644511149
transform -1 0 18032 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1676_
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1677_
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1678_
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1679_
timestamp 1644511149
transform 1 0 10396 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1680_
timestamp 1644511149
transform 1 0 8740 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1681_
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1682_
timestamp 1644511149
transform 1 0 7912 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1683_
timestamp 1644511149
transform 1 0 7728 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1684_
timestamp 1644511149
transform 1 0 7084 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1685_
timestamp 1644511149
transform 1 0 6440 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1686_
timestamp 1644511149
transform 1 0 7728 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1687_
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1688_
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1689_
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1690_
timestamp 1644511149
transform 1 0 17020 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1691_
timestamp 1644511149
transform 1 0 9844 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1692_
timestamp 1644511149
transform 1 0 9476 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1693_
timestamp 1644511149
transform 1 0 12788 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1694_
timestamp 1644511149
transform 1 0 10764 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1695_
timestamp 1644511149
transform 1 0 9108 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1696_
timestamp 1644511149
transform 1 0 10120 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1697_
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1698_
timestamp 1644511149
transform 1 0 9200 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1699_
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1700_
timestamp 1644511149
transform 1 0 10396 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1701_
timestamp 1644511149
transform 1 0 25392 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1702_
timestamp 1644511149
transform 1 0 9384 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1703_
timestamp 1644511149
transform 1 0 9476 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1704_
timestamp 1644511149
transform 1 0 10304 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1705_
timestamp 1644511149
transform 1 0 9660 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1706_
timestamp 1644511149
transform 1 0 10580 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1707_
timestamp 1644511149
transform 1 0 9568 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1708_
timestamp 1644511149
transform 1 0 26036 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1709_
timestamp 1644511149
transform 1 0 14996 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1710_
timestamp 1644511149
transform 1 0 14260 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1711_
timestamp 1644511149
transform 1 0 14812 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1712_
timestamp 1644511149
transform 1 0 13340 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1713_
timestamp 1644511149
transform 1 0 14904 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1714_
timestamp 1644511149
transform 1 0 14720 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1715_
timestamp 1644511149
transform 1 0 14168 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1716_
timestamp 1644511149
transform 1 0 14904 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1717_
timestamp 1644511149
transform 1 0 14904 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1718_
timestamp 1644511149
transform 1 0 15180 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1719_
timestamp 1644511149
transform 1 0 14812 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1720_
timestamp 1644511149
transform 1 0 14444 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1721_
timestamp 1644511149
transform 1 0 17204 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1722_
timestamp 1644511149
transform 1 0 17112 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1723_
timestamp 1644511149
transform 1 0 15916 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1724_
timestamp 1644511149
transform 1 0 16744 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1725_
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1726_
timestamp 1644511149
transform 1 0 15916 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1727_
timestamp 1644511149
transform 1 0 15916 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1728_
timestamp 1644511149
transform 1 0 18400 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1729_
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1730_
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1731_
timestamp 1644511149
transform 1 0 20148 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1732_
timestamp 1644511149
transform 1 0 20976 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1733_
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1734_
timestamp 1644511149
transform 1 0 22080 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1735_
timestamp 1644511149
transform 1 0 22632 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1736_
timestamp 1644511149
transform 1 0 22724 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1737_
timestamp 1644511149
transform 1 0 20240 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1738_
timestamp 1644511149
transform 1 0 17480 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1739_
timestamp 1644511149
transform 1 0 19412 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1740_
timestamp 1644511149
transform 1 0 18032 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _1741_
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1742_
timestamp 1644511149
transform 1 0 16836 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1743_
timestamp 1644511149
transform 1 0 9016 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1744_
timestamp 1644511149
transform 1 0 9752 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1745_
timestamp 1644511149
transform 1 0 12144 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1746_
timestamp 1644511149
transform 1 0 12144 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1747_
timestamp 1644511149
transform 1 0 11316 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1748_
timestamp 1644511149
transform 1 0 10672 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1749_
timestamp 1644511149
transform 1 0 9476 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1750_
timestamp 1644511149
transform 1 0 10028 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1751_
timestamp 1644511149
transform 1 0 8004 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1752_
timestamp 1644511149
transform 1 0 9016 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1753_
timestamp 1644511149
transform 1 0 8188 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1754_
timestamp 1644511149
transform 1 0 7544 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1755_
timestamp 1644511149
transform 1 0 8004 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1756_
timestamp 1644511149
transform 1 0 8464 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _1757_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12420 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1758_
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1759_
timestamp 1644511149
transform 1 0 13156 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1760_
timestamp 1644511149
transform 1 0 15456 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1761_
timestamp 1644511149
transform 1 0 13340 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1762_
timestamp 1644511149
transform 1 0 14720 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1763_
timestamp 1644511149
transform 1 0 13064 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1764_
timestamp 1644511149
transform 1 0 13340 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1765_
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1766_
timestamp 1644511149
transform 1 0 12972 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1767_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1768_
timestamp 1644511149
transform 1 0 11408 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1769_
timestamp 1644511149
transform 1 0 12144 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1770_
timestamp 1644511149
transform 1 0 9384 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1771_
timestamp 1644511149
transform 1 0 7268 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1772_
timestamp 1644511149
transform 1 0 6992 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1773_
timestamp 1644511149
transform 1 0 7728 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1774_
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1775_
timestamp 1644511149
transform 1 0 20700 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1776_
timestamp 1644511149
transform 1 0 17296 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1777_
timestamp 1644511149
transform 1 0 20056 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1778_
timestamp 1644511149
transform 1 0 17296 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1779_
timestamp 1644511149
transform 1 0 21436 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1780_
timestamp 1644511149
transform 1 0 22540 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1781_
timestamp 1644511149
transform 1 0 23552 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1782_
timestamp 1644511149
transform 1 0 11684 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1783_
timestamp 1644511149
transform 1 0 14352 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1784_
timestamp 1644511149
transform 1 0 16928 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1785_
timestamp 1644511149
transform 1 0 15456 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dlxtn_1  _1786_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23460 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1787_
timestamp 1644511149
transform 1 0 24932 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1788_
timestamp 1644511149
transform 1 0 22724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1789_
timestamp 1644511149
transform 1 0 19872 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1790_
timestamp 1644511149
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1791_
timestamp 1644511149
transform 1 0 20976 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1792_
timestamp 1644511149
transform 1 0 21988 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1793_
timestamp 1644511149
transform 1 0 21896 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1794_
timestamp 1644511149
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  _1795_
timestamp 1644511149
transform 1 0 15548 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1796_
timestamp 1644511149
transform 1 0 9568 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1797_
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1798_
timestamp 1644511149
transform 1 0 6992 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1799_
timestamp 1644511149
transform 1 0 6808 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1800_
timestamp 1644511149
transform 1 0 6992 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1801_
timestamp 1644511149
transform 1 0 8004 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1802_
timestamp 1644511149
transform 1 0 9568 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1803_
timestamp 1644511149
transform 1 0 10764 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dlxtn_1  _1804_
timestamp 1644511149
transform 1 0 18584 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1805_
timestamp 1644511149
transform 1 0 19320 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1806_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17112 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtp_1  _1807_
timestamp 1644511149
transform 1 0 17664 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1808_
timestamp 1644511149
transform 1 0 17664 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1809_
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1810_
timestamp 1644511149
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1811_
timestamp 1644511149
transform 1 0 21528 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1812_
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1813_
timestamp 1644511149
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1814_
timestamp 1644511149
transform 1 0 18124 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1815_
timestamp 1644511149
transform 1 0 20700 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1816_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25116 0 1 16320
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1817_
timestamp 1644511149
transform 1 0 9844 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dlxtn_1  _1818_
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1819_
timestamp 1644511149
transform 1 0 21988 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1820_
timestamp 1644511149
transform 1 0 20240 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_2  _1821_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20424 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_1  _1822_
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1823_
timestamp 1644511149
transform 1 0 18308 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1824_
timestamp 1644511149
transform 1 0 19596 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1825_
timestamp 1644511149
transform 1 0 16836 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1826_
timestamp 1644511149
transform 1 0 20976 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1827_
timestamp 1644511149
transform 1 0 16376 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1828_
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1829_
timestamp 1644511149
transform 1 0 15088 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1830_
timestamp 1644511149
transform 1 0 14444 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1831_
timestamp 1644511149
transform 1 0 14352 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_1  _1832_
timestamp 1644511149
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__dlxtn_2  _1833_
timestamp 1644511149
transform 1 0 14168 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__dlxtn_1  _1834_
timestamp 1644511149
transform 1 0 15732 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_2  _1835_
timestamp 1644511149
transform 1 0 25944 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1836_
timestamp 1644511149
transform 1 0 14352 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1837_
timestamp 1644511149
transform 1 0 14444 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1838_
timestamp 1644511149
transform 1 0 14168 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1839_
timestamp 1644511149
transform 1 0 14444 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1840_
timestamp 1644511149
transform 1 0 14996 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1841_
timestamp 1644511149
transform 1 0 17204 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1842_
timestamp 1644511149
transform 1 0 14720 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1843_
timestamp 1644511149
transform 1 0 15640 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1844_
timestamp 1644511149
transform 1 0 17664 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1845_
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1846_
timestamp 1644511149
transform 1 0 19872 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1847_
timestamp 1644511149
transform 1 0 21620 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1848_
timestamp 1644511149
transform 1 0 22172 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1849_
timestamp 1644511149
transform 1 0 16744 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1850_
timestamp 1644511149
transform 1 0 9476 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1851_
timestamp 1644511149
transform 1 0 10948 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1852_
timestamp 1644511149
transform 1 0 11684 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1853_
timestamp 1644511149
transform 1 0 10304 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1854_
timestamp 1644511149
transform 1 0 8188 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1855_
timestamp 1644511149
transform 1 0 7176 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1856_
timestamp 1644511149
transform 1 0 6992 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1857_
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19688 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_clk
timestamp 1644511149
transform 1 0 17848 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_clk
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1
timestamp 1644511149
transform 1 0 30728 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1644511149
transform 1 0 23552 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input4
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1644511149
transform 1 0 10396 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1644511149
transform 1 0 37812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1644511149
transform 1 0 37812 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1644511149
transform 1 0 20700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1644511149
transform 1 0 37812 0 -1 13056
box -38 -48 406 592
<< labels >>
rlabel metal5 s 1104 20616 38824 20936 6 VGND
port 0 nsew ground input
rlabel metal4 s 19568 2128 19888 37584 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 5298 38824 5618 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 35934 38824 36254 6 VPWR
port 1 nsew power input
rlabel metal4 s 4208 2128 4528 37584 6 VPWR
port 1 nsew power input
rlabel metal4 s 34928 2128 35248 37584 6 VPWR
port 1 nsew power input
rlabel metal3 s 39200 23128 40000 23248 6 clk
port 2 nsew signal input
rlabel metal2 s 13542 39200 13598 40000 6 led_flag
port 3 nsew signal tristate
rlabel metal2 s 30930 0 30986 800 6 restart
port 4 nsew signal input
rlabel metal2 s 23846 39200 23902 40000 6 rotary_a
port 5 nsew signal input
rlabel metal2 s 18 0 74 800 6 rotary_b
port 6 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 rst
port 7 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 select
port 8 nsew signal input
rlabel metal3 s 39200 1368 40000 1488 6 seven_segment_digit
port 9 nsew signal tristate
rlabel metal3 s 0 10888 800 11008 6 seven_segment_out[0]
port 10 nsew signal tristate
rlabel metal3 s 39200 34008 40000 34128 6 seven_segment_out[1]
port 11 nsew signal tristate
rlabel metal2 s 34150 39200 34206 40000 6 seven_segment_out[2]
port 12 nsew signal tristate
rlabel metal2 s 20626 0 20682 800 6 seven_segment_out[3]
port 13 nsew signal tristate
rlabel metal3 s 0 32648 800 32768 6 seven_segment_out[4]
port 14 nsew signal tristate
rlabel metal2 s 3238 39200 3294 40000 6 seven_segment_out[5]
port 15 nsew signal tristate
rlabel metal3 s 39200 12248 40000 12368 6 seven_segment_out[6]
port 16 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
